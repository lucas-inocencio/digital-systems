-- ALU 4-bit

-- The operations to be performed in the ALU must be selected by control inputs.
-- work must have 3 external switches (switchers) to control such operations.
-- Mandatory operations: addition, subtraction in 2's complement, increment +1, exchange of signal.
-- Students will have to develop an auxiliary module that will be used to vary the operands input that will test the ALU.
-- The input data and the result of the operation must be displayed on the LEDs available on the FPGA board.
-- ALU outputs must be the result and the four flags (Zero, negative, carry out, overflow) which should be shown on the LEDs. Operation:
-- The input operands are generated by an auxiliary module that will contain a contactor that
-- will loop through all binaries represented by 4 bits. Entries are shown simultaneously
-- in the LEDs. Then, the ALU receives the operands and produces the result also shown in the
-- 7 segment display. Furthermore, the ALU generates 4 flags that are shown on the LEDs.
-- The ALU inputs are generated by an auxiliary module, a counter, part
-- member of the project. The two entries are shown, together with the result, in the
-- 7-segment displays available. The LEDs are used to show the four “flags”. You
-- operands change, in ascending order, every 2 seconds.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ALU is
    Port ( A, B : in  STD_LOGIC_VECTOR (3 downto 0);
           Selector : in  STD_LOGIC_VECTOR (2 downto 0);
           Flags : out  STD_LOGIC_VECTOR (3 downto 0);
           ALU_Output : out  STD_LOGIC_VECTOR (3 downto 0));
end ALU;

architecture Behavioral of ALU is

begin

process(A, B, Selector)
begin
    case Selector is
        when "000" => ALU_Output <= A + B; -- Addition
        when "001" => ALU_Output <= A - B; -- Subtraction in 2's complement
        when "010" => ALU_Output <= A + 1; -- Increment +1
        when "011" => ALU_Output <= B; -- Exchange of signal
        when "100" => ALU_Output <= A and B; -- AND
        when "101" => ALU_Output <= A or B; -- OR
        when "110" => ALU_Output <= A xor B; -- XOR
        when "111" => ALU_Output <= A nand B; -- NAND
        when others => ALU_Output <= "0000";
    end case;
end process;

process(ALU_Output)
begin
    if ALU_Output = "0000" then
        Flags <= "1000";
    elsif ALU_Output < "0000" then
        Flags <= "0100";
    elsif ALU_Output > "1111" then
        Flags <= "0010";
    else
        Flags <= "0001";
    end if;
end process;

end Behavioral;