// ALU