From: <Saved by Blink>
Snapshot-Content-Location: https://drive.google.com/file/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view
Subject: decoder7seg.vhd - Google Drive
Date: Tue, 20 Jun 2023 16:36:22 -0000
MIME-Version: 1.0
Content-Type: multipart/related;
	type="text/html";
	boundary="----MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----"


------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/html
Content-ID: <frame-419165DDFD6EFAABF68E51E9196DF57B@mhtml.blink>
Content-Transfer-Encoding: binary
Content-Location: https://drive.google.com/file/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view

<!DOCTYPE html><html><head><meta http-equiv="Content-Type" content="text/html; charset=UTF-8"><link rel="stylesheet" type="text/css" href="cid:css-62abb5c1-8626-4e4f-95af-4454145f1290@mhtml.blink" /><link rel="stylesheet" type="text/css" href="cid:css-d28e6a9c-e182-4cb7-87e1-14d2709c3aca@mhtml.blink" /><meta name="google" content="notranslate"><meta http-equiv="X-UA-Compatible" content="IE=edge;"><meta name="viewport" content="width=device-width, initial-scale=1.0, maximum-scale=1.0, minimum-scale=1.0, user-scalable=0"><meta name="referrer" content="origin"><title>decoder7seg.vhd - Google Drive</title><meta property="og:title" content="decoder7seg.vhd"><meta property="og:type" content="article"><meta property="og:site_name" content="Google Docs"><meta property="og:url" content="https://drive.google.com/file/u/0/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view?usp=drive_web&amp;usp=embed_facebook"><link rel="shortcut icon" href="https://ssl.gstatic.com/images/branding/product/1x/drive_2020q4_32dp.png"><link rel="stylesheet" href="https://fonts.googleapis.com/css?family=Google+Sans_old:300,400,500,700" nonce=""><link rel="stylesheet" href="https://www.gstatic.com/_/apps-fileview/_/ss/k=apps-fileview.v.omJv0zZNxLk.L.W.O/am=AAAE/d=0/rs=AO0039tfU3F6Yks5o2y0ftEU4qi8duRDBA" nonce=""><link type="text/css" rel="stylesheet" href="https://www.gstatic.com/og/_/ss/k=og.qtm.Bcf36HdLxAc.L.W.O/m=qcwid/excm=qaaw,qadd,qaid,qein,qhaw,qhba,qhbr,qhch,qhga,qhid,qhin/d=1/ed=1/ct=zgms/rs=AA2YrTtrdJEPAVAbPPca5uf3TCfVu9JrgA" nonce=""></head><body dir="ltr" role="application" itemscope="" itemtype="http://schema.org/CreativeWork/FileObject" class="ndfHFb-c4YZDc-uoC0bf ndfHFb-c4YZDc-qbOKL-OEVmcd" jsaction="UjQMac:.CLIENT"><div style="display:none" aria-hidden="true"><div id="one-google-bar" class="ndfHFb-c4YZDc-Woal0c-jcJzye-ZMv3u ndfHFb-c4YZDc-n1UuX-Bz112c"><div class="gb_Pa gb_f gb_gb gb_i gb_Rc gb_Ha gb_Qa" id="gb" style="background-color:transparent"><div class="gb_Dd gb_eb gb_sd" ng-non-bindable="" data-ogsr-up="" style="padding:0;height:auto;display:block"><div class="gb_Xd" style="display:block"><div class="gb_9c"></div><div class="gb_b gb_Rd gb_3f gb_x gb_Pb gb_Ud"><div class="gb_g gb_db gb_3f gb_x"><a class="gb_d gb_Fa gb_x" aria-label="Conta do Google: Roberto Gonçalves Pacheco  
(robertopacheco@poli.ufrj.br)" href="https://accounts.google.com/SignOutOptions?hl=pt-BR&amp;continue=https://drive.google.com/file/u/0/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view%3Fusp%3Ddrive_web&amp;service=writely&amp;ec=GBRAGQ" role="button" tabindex="0"><img class="gb_k gbii" src="https://lh3.googleusercontent.com/ogw/AOLn63Fd7vZE5o2FaKK7Sg0PDYjfXo_g8YLZTYOwvcVc=s32-c-mo" alt="" aria-hidden="true" data-noaft=""></a><div class="gb_jb"></div><div class="gb_ib"></div></div></div></div><div style="overflow: hidden; position: absolute; top: 0px; visibility: hidden; width: 400px; z-index: 991; height: 0px; margin-top: 57px; right: 0px; margin-right: 4px;"></div></div></div></div></div><meta itemprop="name" content="decoder7seg.vhd" aria-hidden="true"><meta itemprop="faviconUrl" content="https://ssl.gstatic.com/images/branding/product/1x/drive_2020q4_32dp.png" aria-hidden="true"><meta itemprop="url" content="https://drive.google.com/file/u/0/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view?usp=drive_web&amp;usp=embed_googleplus" aria-hidden="true"><div ng-non-bindable="" aria-hidden="true"></div><div class="gb_n" ng-non-bindable="" aria-hidden="true"><div class="gb_Ic"><div>Conta do Google</div><div class="gb_Hb">Roberto Gonçalves Pacheco</div><div>robertopacheco@poli.ufrj.br</div></div></div><div class="ndfHFb-c4YZDc ndfHFb-c4YZDc-AHmuwe-Hr88gd-OWB6Me dif24c vhoiae LgGVmb bvmRsc ndfHFb-c4YZDc-N4imRe ndfHFb-c4YZDc-vyDMJf-aZ2wEe ndfHFb-c4YZDc-i5oIFb ndfHFb-c4YZDc-uoC0bf ndfHFb-c4YZDc-TSZdd" aria-label="Mostrando leitor." tabindex="0"><div class="ndfHFb-c4YZDc-bnBfGc ndfHFb-c4YZDc-zTETae" tabindex="0" aria-label="Nenhuma visualização disponível"></div><div class="ndfHFb-c4YZDc-JNEHMb"><div class="ndfHFb-c4YZDc-uWtm3-ORHb" role="status" tabindex="0"><div class="ndfHFb-c4YZDc-uWtm3-ORHb-Bz112c"></div><div class="ndfHFb-c4YZDc-uWtm3-ORHb-bN97Pc"><div class="ndfHFb-c4YZDc-uWtm3-ORHb-Ne3sFf"></div><div class="ndfHFb-c4YZDc-uWtm3-ORHb-LQLjdd"><div class="ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Pedir análise</div></div><div class="ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Saiba mais</div></div><div class="ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe" title="" role="button" aria-label="Dispensar aviso" tabindex="0" style="user-select: none;"><div class="ndfHFb-c4YZDc-Bz112c  ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-Bz112c" aria-label="Fechar banner"></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf"><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Bz112c"></div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-bN97Pc"><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-jOfkMb">Assinatura pendente</div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Vkfede-Ne3sFf"></div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-LQLjdd"><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Assinar</div></div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Rejeitar</div></div><div class="ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Ver detalhes</div></div></div></div></div><div class="ndfHFb-c4YZDc-L7w45e-ORHb" role="status" tabindex="0"><div class="ndfHFb-c4YZDc-L7w45e-ORHb-Bz112c"></div><div class="ndfHFb-c4YZDc-L7w45e-ORHb-bN97Pc"><div class="ndfHFb-c4YZDc-L7w45e-ORHb-Ne3sFf"></div><div class="ndfHFb-c4YZDc-L7w45e-ORHb-LQLjdd"><div class="ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Não é spam</div></div><div class="ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Remover permanentemente</div></div><div class="ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe" title="" role="button" aria-label="Dispensar aviso" tabindex="0" style="user-select: none;"><div class="ndfHFb-c4YZDc-Bz112c  ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-Bz112c" aria-label="Fechar banner"></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb" role="status" tabindex="0"><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Bz112c"></div><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-bN97Pc"><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Ne3sFf"></div><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-LQLjdd"><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe" title="" role="button" tabindex="0" style="user-select: none;">Não é spam</div></div><div class="ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-LgbsSe-sM5MNb"><div class="VIpgJd-TzA9Ye-eEGnhe VIpgJd-C41vtd-LgbsSe" title="" role="button" aria-label="Dispensar aviso" tabindex="0" style="user-select: none;"><div class="ndfHFb-c4YZDc-Bz112c  ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c" aria-label="Fechar banner"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-K9a4Re" style="bottom: 0px; top: 0px;"><div class="ndfHFb-c4YZDc-E7ORLb-LgbsSe ndfHFb-c4YZDc-LgbsSe-OWB6Me ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e" role="button" aria-disabled="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="r,c" data-tooltip-offset="-6" style="user-select: none; left: 16px; display: none;"><div class="ndfHFb-c4YZDc-DH6Rkf-AHe6Kc"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-tJiF1e-LgbsSe ndfHFb-c4YZDc-LgbsSe-OWB6Me ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e" role="button" aria-disabled="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="l,c" data-tooltip-offset="-6" style="user-select: none; right: 16px; display: none;"><div class="ndfHFb-c4YZDc-DH6Rkf-AHe6Kc"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-q77wGc ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e"><div class="ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb" style="display: none;"></div><div class="ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb" style="display: none;"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-m9bMae-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Diminuir o zoom" data-tooltip="Diminuir o zoom" style="user-select: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe VIpgJd-TzA9Ye-eEGnhe" role="button" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" style="user-select: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-bEDTcc-LgbsSe VIpgJd-TzA9Ye-eEGnhe" role="button" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" style="user-select: none;" aria-label="Aumentar o zoom" data-tooltip="Aumentar o zoom"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-LzGo7c" style="display: none;"></div></div><div class="ndfHFb-c4YZDc-K9a4Re-nKQ6qf ndfHFb-c4YZDc-TvD9Pc-qnnXGd" role="main" style=""><div class="ndfHFb-c4YZDc-EglORb-ge6pde ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf" role="status" tabindex="-1" aria-label="Carregando" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div><span class="ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" aria-hidden="true">Carregando…</span></div><div style="display:none" id="drive-active-item-info">{"id": "1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3", "title": "decoder7seg.vhd", "mimeType": "application\/x-virtualbox-vhd"}</div><div style="display: none;"></div><div class="ndfHFb-c4YZDc-EglORb-u0pjoe ndfHFb-c4YZDc-neVct-RCfa3e" style="left: 12px; top: 64px;"><div class="ndfHFb-c4YZDc-EglORb-haAclf ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" tabindex="-1"><div class="ndfHFb-c4YZDc-EglORb-u0pjoe-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" tabindex="-1">Nenhuma visualização disponível</div><div class="ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf" style="display: none;"><a class="ndfHFb-c4YZDc-EglORb-u0pjoe-KY1xSc-z5C9Gb-hSRGPd" href="https://drive.google.com/file/d/1xFe4zzI8xE2AY5OmdpEHGZSbnjZqGAn3/view">Saiba mais</a></div><div class="ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" tabindex="-1" style="display: none;"></div><pre class="ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" tabindex="-1" style="display: none;"></pre><div class="ndfHFb-c4YZDc-EglORb-joDrKf-u0pjoe-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" style="display: none;">Tentando novamente…</div><div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe" role="button" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Fazer o download" data-tooltip="Fazer o download"><div class="ndfHFb-c4YZDc-nupQLb-Bz112c ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-Bz112c"></div><div class="ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-fmcmS" aria-hidden="true">Download</div></div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe" style="display: none;"><div class="ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-Bz112c"></div><div class="ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-fmcmS">Conectar mais apps…</div></div></div></div><div class="ndfHFb-c4YZDc-rovI0b-haAclf" style="display: none;"></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e" role="toolbar"><div class="ndfHFb-c4YZDc-Wrql6b-SmKAyb" style="margin-right: 12px; padding-left: 12px;"><div class="ndfHFb-c4YZDc-Wrql6b-hOcTPc" style="left: 12px;"><div class="ndfHFb-c4YZDc-Wrql6b-Bz112c" tabindex="-1" role="img" aria-label="Ícone de Arquivo desconhecido" style="background-image: url(&quot;https://drive-thirdparty.googleusercontent.com/32/type/application/x-virtualbox-vhd&quot;); background-position: left top; background-repeat: no-repeat;"></div><div class="ndfHFb-c4YZDc-Wrql6b-jfdpUb" tabindex="-1"><div class="ndfHFb-c4YZDc-Wrql6b-V1ur5d" aria-label="decoder7seg.vhd" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip="decoder7seg.vhd"> ... </div><div class="ndfHFb-c4YZDc-Wrql6b-V1ur5d ndfHFb-c4YZDc-Wrql6b-V1ur5d-hpYHOb">d ... d</div><div class="ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d" style="display: none;"></div><div class="ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-hpYHOb"></div></div><div class="ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c" style="display: none;"></div><div class="ndfHFb-c4YZDc-TL3Ynd-V67aGc-haAclf ndfHFb-c4YZDc-LgbsSe-OWB6Me" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-disabled="true"></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-C7uZwb-ibnC6b-Btuy5e ndfHFb-c4YZDc-LgbsSe-OWB6Me" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-disabled="true" aria-hidden="true" aria-label="Bloqueado" data-tooltip="Bloqueado" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c ndfHFb-c4YZDc-pGuBYc-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-DdWCyb-b0t70b" style="display: none;"><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d" style="display: none;"><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c" style="display: none;"></div><div class="ndfHFb-c4YZDc-FNFY6c-V67aGc">Abrir</div></div><div class="ndfHFb-c4YZDc-Wrql6b-PlOyMe ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" style="user-select: none; display: none;" aria-hidden="true"><div class="ndfHFb-c4YZDc-Wrql6b-PlOyMe-bN97Pc">Extrair</div><div class="ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" aria-expanded="false" aria-haspopup="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Abrir com" data-tooltip="Abrir com" style="user-select: none; display: none;" aria-hidden="true"><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe"></div><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb"><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS" tabindex="-1">Abrir com</div><div class="ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b" style="display: none;"><div class="ndfHFb-c4YZDc-zM6fo-GMvhG-Bz112c ndfHFb-c4YZDc-Bz112c"></div><span class="ndfHFb-c4YZDc-zM6fo-GMvhG-fmcmS" tabindex="0" role="alert"></span></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b"><div class="ndfHFb-c4YZDc-GSQQnc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe" aria-label="Ver em outra janela" style="display: none;"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-LQLjdd"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb" style="display: none;"><div><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c ndfHFb-c4YZDc-LgbsSe-OWB6Me" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-disabled="true" aria-hidden="true" aria-label="Fazer o download" data-tooltip="Fazer o download" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c ndfHFb-c4YZDc-nupQLb-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-z5C9Gb-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" aria-expanded="false" aria-haspopup="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Mais ações" data-tooltip="Mais ações" style="user-select: none;" aria-hidden="false" tabindex="0"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div></div><div class="ndfHFb-c4YZDc-n1UuX-Bz112c" title="Roberto Gonçalves Pacheco 
(robertopacheco@poli.ufrj.br)"><img src="https://lh3.googleusercontent.com/a/AAcHTtdQDe6r_XGCNEiOx6KZzpjviLw9RqZeAy_GGnpv=s50-c-k-no" class="ndfHFb-c4YZDc-n1UuX-RJLb9c" alt="Roberto Gonçalves Pacheco 
(robertopacheco@poli.ufrj.br)" tabindex="0"></div></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-b0t70b ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce" aria-hidden="true"><div class="ndfHFb-c4YZDc-MZArnb-b0t70b-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-tJHJj"><div class="ndfHFb-c4YZDc-MZArnb-cXCLoc ndfHFb-c4YZDc-MZArnb-cXCLoc-DKlKme ndfHFb-c4YZDc-MZArnb-cXCLoc-ma6Yeb" role="tablist" aria-label="Barra de guias do painel de detalhes. Pressione as teclas de seta esquerda e direita para mudar de guia." aria-activedescendant="dvdt_goog_508823002" style="user-select: none;"><div class="ndfHFb-c4YZDc-MZArnb-AznF2e ndfHFb-c4YZDc-MZArnb-AznF2e-ZmdkE ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd" role="tab" aria-selected="true" id="dvdt_goog_508823002" tabindex="0" style="user-select: none;">Detalhes</div><div class="ndfHFb-c4YZDc-MZArnb-AznF2e ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge" role="tab" aria-selected="false" id="dvdt_goog_508823003" style="user-select: none; display: none;" aria-hidden="true">Comentários</div></div><div class="ndfHFb-c4YZDc-TvD9Pc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" style="user-select: none;" aria-label="Ocultar detalhes" data-tooltip="Ocultar detalhes"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-bN97Pc ndfHFb-c4YZDc-s2gQvd"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-nUpftc" role="tabpanel" aria-labelledby="dvdt_goog_508823002" style=""><div role="complementary" aria-label="Informações gerais" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Informações gerais</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Tipo</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">Arquivo desconhecido</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Dimensões</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Tamanho</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">820 bytes</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Duração</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Local</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"><div class="ndfHFb-c4YZDc-MZArnb-P86uke-PntVL"><div><div class="ndfHFb-c4YZDc-MZArnb-P86uke-Bz112c" style="background-image: url(https://drive-thirdparty.googleusercontent.com/16/type/application/vnd.google-apps.folder+shared); background-size:cover;"></div><div class="ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd ndfHFb-c4YZDc-LgbsSe" role="button" tabindex="0" data-id="19zi4nQFPgWUFUtTY9vwwX9hh24FaGoqlMGddVXd2xIqd2VKyYKp1jp8uh-KUOuOyhNP0J1R3" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip="Sistemas Digitais 2022-2" data-tooltip-only-on-overflow="true" style="user-select: none;">Sistemas Digitais 2022-2</div></div></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Modificado</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">13:36 12 de out. de 2022</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Criado</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">13:37 12 de out. de 2022</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Aberto por mim</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">13:37 12 de out. de 2022</div></div></div></div></div><div role="complementary" aria-label="Compartilhamento" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Compartilhamento</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-BA389-V67aGc"><div class="ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c"><div class="ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e" data-tooltip="Sistemas_Digitais_2022_2_teachers_c3fff74d@poli.ufrj.br" aria-label="Sistemas_Digitais_2022_2_teachers_c3fff74d@poli.ufrj.br" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-MZArnb-YLEF4c-Bz112c ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c" role="img" alt=""></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d" data-tooltip="Professores de Sistemas Digitais 2022-2" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip-only-on-overflow="true">Professores de Sistemas Digitais 2022-2</div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-nNAX0">Pode editar</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-BA389-V67aGc"><div class="ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c"><div class="ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e" data-tooltip="Sistemas_Digitais_2022_2_39aaa311@poli.ufrj.br" aria-label="Sistemas_Digitais_2022_2_39aaa311@poli.ufrj.br" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-MZArnb-YLEF4c-Bz112c ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c" role="img" alt=""></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d" data-tooltip="Sistemas Digitais 2022-2" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip-only-on-overflow="true">Sistemas Digitais 2022-2</div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-nNAX0">Pode ver</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-BA389-V67aGc"><div class="ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c"><img class="ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c" alt="" src="https://lh3.googleusercontent.com/a/AAcHTtdQDe6r_XGCNEiOx6KZzpjviLw9RqZeAy_GGnpv=s64" role="img" data-tooltip="robertopacheco@poli.ufrj.br" aria-label="robertopacheco@poli.ufrj.br" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6"></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d" data-tooltip="Roberto Gonçalves Pacheco" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip-only-on-overflow="true">Roberto Gonçalves Pacheco</div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-nNAX0">Proprietário</div></div></div></div></div><div role="complementary" aria-label="Descrição" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Descrição</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" aria-label="Editar a descrição" data-tooltip="Editar a descrição" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div><div class="ndfHFb-c4YZDc-MZArnb-ij8cu" role="complementary" tabindex="0">Nenhuma descrição</div><textarea class="ndfHFb-c4YZDc-MZArnb-ij8cu-DyVDA ndfHFb-c4YZDc-s2gQvd" role="textbox" aria-multiline="true" style="display: none;"></textarea></div></div></div><div role="complementary" aria-label="Permissão para download" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Permissão para download</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" style="user-select: none; display: none;"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-nupQLb-BA389-Ne3sFf" id="dvddp_goog_508823001">Os leitores podem fazer o download</div></div></div></div><div></div></div><div class="ndfHFb-c4YZDc-MZArnb-RDNXzf-nUpftc" role="tabpanel" aria-labelledby="dvdt_goog_508823003" style="display: none;"></div></div></div></div><div class="VIpgJd-TUo6Hb-xJ5Hnf ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-xJ5Hnf" style="display: none;"></div><div class="VIpgJd-TUo6Hb ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-haAclf" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe" role="status" tabindex="-1" aria-label="Carregando" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div><span class="ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" aria-hidden="true">Carregando…</span></div></div><span tabindex="0" style="display: none; position: absolute;"></span><div class="ndfHFb-c4YZDc-zsEIvc-b0t70b ndfHFb-c4YZDc-zsEIvc-MqcBrc-b0t70b" style="display: none; top: 64px;"></div></div><span class="ndfHFb-c4YZDc-AznF2e-DTMEae" tabindex="0" style="" aria-hidden="true"></span><iframe id="apiproxy82411c4c82d95adef5e7dae7c39b0f518a351d020.2872649575" name="apiproxy82411c4c82d95adef5e7dae7c39b0f518a351d020.2872649575" src="cid:frame-8DF312FC58F6EE99A3ED96B5411FF620@mhtml.blink" tabindex="-1" aria-hidden="true" style="width: 1px; height: 1px; position: absolute; top: -100px; display: none;"></iframe><div id="goog-lr-9" aria-live="polite" aria-atomic="true" style="position: absolute; top: -1000px; height: 1px; overflow: hidden;">Nenhuma visualização disponível</div></body></html>
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/css
Content-Transfer-Encoding: binary
Content-Location: cid:css-62abb5c1-8626-4e4f-95af-4454145f1290@mhtml.blink

@charset "utf-8";

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xFIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+460-52F, U+1C80-1C88, U+20B4, U+2DE0-2DFF, U+A640-A69F, U+FE2E-FE2F; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xMIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xEIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+1F00-1FFF; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xLIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xHIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xGIzIXKMnyrYk.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: Roboto; font-style: italic; font-weight: 400; src: local("Roboto Italic"), local("Roboto-Italic"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOkCnqEu92Fr1Mu51xIIzIXKMny.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fCRc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+460-52F, U+1C80-1C88, U+20B4, U+2DE0-2DFF, U+A640-A69F, U+FE2E-FE2F; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fABc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fCBc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+1F00-1FFF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fBxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fCxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fChc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 300; src: local("Roboto Light"), local("Roboto-Light"), local("sans-serif-light"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmSU5fBBc4AMP6lQ.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu72xKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+460-52F, U+1C80-1C88, U+20B4, U+2DE0-2DFF, U+A640-A69F, U+FE2E-FE2F; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu5mxKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7mxKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+1F00-1FFF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu4WxKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7WxKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7GxKKTU1Kvnz.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 400; src: local("Roboto Regular"), local("Roboto-Regular"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu4mxKKTU1Kg.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCRc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+460-52F, U+1C80-1C88, U+20B4, U+2DE0-2DFF, U+A640-A69F, U+FE2E-FE2F; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fABc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCBc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+1F00-1FFF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fBxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fChc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 500; src: local("Roboto Medium"), local("Roboto-Medium"), local("sans-serif-medium"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fBBc4AMP6lQ.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCRc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+460-52F, U+1C80-1C88, U+20B4, U+2DE0-2DFF, U+A640-A69F, U+FE2E-FE2F; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfABc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCBc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+1F00-1FFF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfBxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCxc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfChc4AMP6lbBP.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: Roboto; font-style: normal; font-weight: 700; src: local("Roboto Bold"), local("Roboto-Bold"), local("sans-serif"), url("//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfBBc4AMP6lQ.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/css
Content-Transfer-Encoding: binary
Content-Location: cid:css-d28e6a9c-e182-4cb7-87e1-14d2709c3aca@mhtml.blink

@charset "utf-8";

.gb_gb:not(.gb_ld) { font: 13px / 27px Roboto, Arial, sans-serif; z-index: 986; }

@-webkit-keyframes gb__a { 
  0% { opacity: 0; }
  50% { opacity: 1; }
}

@keyframes gb__a { 
  0% { opacity: 0; }
  50% { opacity: 1; }
}

a.gb_ka { border: none; color: rgb(66, 133, 244); cursor: default; font-weight: bold; outline: none; position: relative; text-align: center; text-decoration: none; text-transform: uppercase; white-space: nowrap; user-select: none; }

a.gb_ka:hover::after, a.gb_ka:focus::after { background-color: rgba(0, 0, 0, 0.12); content: ""; height: 100%; left: 0px; position: absolute; top: 0px; width: 100%; }

a.gb_ka:hover, a.gb_ka:focus { text-decoration: none; }

a.gb_ka:active { background-color: rgba(153, 153, 153, 0.4); text-decoration: none; }

a.gb_la { background-color: rgb(66, 133, 244); color: rgb(255, 255, 255); }

a.gb_la:active { background-color: rgb(0, 67, 178); }

.gb_ma { box-shadow: rgba(0, 0, 0, 0.16) 0px 1px 1px; }

.gb_ka, .gb_la, .gb_na, .gb_oa { display: inline-block; line-height: 28px; padding: 0px 12px; border-radius: 2px; }

.gb_na { background: rgb(248, 248, 248); border: 1px solid rgb(198, 198, 198); }

.gb_oa { background: rgb(248, 248, 248); }

.gb_na, #gb a.gb_na.gb_na, .gb_oa { color: rgb(102, 102, 102); cursor: default; text-decoration: none; }

#gb a.gb_oa { cursor: default; text-decoration: none; }

.gb_oa { border: 1px solid rgb(66, 133, 244); font-weight: bold; outline: none; background: -webkit-linear-gradient(top, rgb(67, 135, 253), rgb(70, 131, 234)); }

#gb a.gb_oa { color: rgb(255, 255, 255); }

.gb_oa:hover { box-shadow: rgba(0, 0, 0, 0.15) 0px 1px 0px; }

.gb_oa:active { box-shadow: rgba(0, 0, 0, 0.15) 0px 2px 0px inset; background: -webkit-linear-gradient(top, rgb(60, 122, 228), rgb(63, 118, 211)); }

#gb .gb_pa { background: rgb(255, 255, 255); border: 1px solid rgb(218, 220, 224); color: rgb(26, 115, 232); display: inline-block; text-decoration: none; }

#gb .gb_pa:hover { background: rgb(248, 251, 255); border-color: rgb(218, 220, 224); color: rgb(23, 78, 166); }

#gb .gb_pa:focus { background: rgb(244, 248, 255); color: rgb(23, 78, 166); outline: rgb(23, 78, 166) solid 1px; }

#gb .gb_pa:active, #gb .gb_pa:focus:active { background: rgb(236, 243, 254); color: rgb(23, 78, 166); }

#gb .gb_pa.gb_i { background: transparent; border: 1px solid rgb(95, 99, 104); color: rgb(138, 180, 248); text-decoration: none; }

#gb .gb_pa.gb_i:hover { background: rgba(255, 255, 255, 0.04); color: rgb(232, 234, 237); }

#gb .gb_pa.gb_i:focus { background: rgba(232, 234, 237, 0.12); color: rgb(232, 234, 237); outline: rgb(232, 234, 237) solid 1px; }

#gb .gb_pa.gb_i:active, #gb .gb_pa.gb_i:focus:active { background: rgba(232, 234, 237, 0.1); color: rgb(232, 234, 237); }

.gb_m { display: none !important; }

.gb_1a { visibility: hidden; }

.gb_Rd { display: inline-block; vertical-align: middle; }

.gb_Td .gb_l { bottom: -3px; right: -5px; }

.gb_g { position: relative; }

.gb_d { display: inline-block; outline: none; vertical-align: middle; border-radius: 2px; box-sizing: border-box; height: 40px; width: 40px; cursor: pointer; text-decoration: none; }

#gb#gb a.gb_d { cursor: pointer; text-decoration: none; }

.gb_d, a.gb_d { color: rgb(0, 0, 0); }

.gb_ib { border-color: transparent transparent rgb(255, 255, 255); border-style: dashed dashed solid; border-width: 0px 8.5px 8.5px; display: none; position: absolute; left: 11.5px; top: 33px; z-index: 1; height: 0px; width: 0px; animation: 0.2s ease 0s 1 normal none running gb__a; }

.gb_jb { border-color: transparent transparent rgba(0, 0, 0, 0.2); border-style: dashed dashed solid; border-width: 0px 8.5px 8.5px; display: none; position: absolute; left: 11.5px; z-index: 1; height: 0px; width: 0px; animation: 0.2s ease 0s 1 normal none running gb__a; top: 32px; }

.gb_U { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.2); color: rgb(0, 0, 0); box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 10px; display: none; outline: none; overflow: hidden; position: absolute; right: 8px; top: 62px; animation: 0.2s ease 0s 1 normal none running gb__a; border-radius: 2px; user-select: text; }

.gb_Rd.gb_La .gb_ib, .gb_Rd.gb_La .gb_jb, .gb_Rd.gb_La .gb_U, .gb_La.gb_U { display: block; }

.gb_Rd.gb_La.gb_Ud .gb_ib, .gb_Rd.gb_La.gb_Ud .gb_jb { display: none; }

.gb_Vd { position: absolute; right: 8px; top: 62px; z-index: -1; }

.gb_7a .gb_ib, .gb_7a .gb_jb, .gb_7a .gb_U { margin-top: -10px; }

.gb_Rd:first-child, #gbsfw:first-child + .gb_Rd { padding-left: 4px; }

.gb_Pa.gb_Wd .gb_Rd:first-child { padding-left: 0px; }

.gb_Xd { position: relative; }

.gb_Pa .gb_Zd .gb_Pd.gb_od, .gb_Pa.gb_Qa .gb_Zd .gb_Pd.gb_od { padding: 3px 8px 3px 16px; }

.gb_Zd .gb_0d { display: inline-block; }

.gb_Zd .gb_od { border-radius: 100px; background: rgb(11, 87, 208); color: rgb(255, 255, 255); font-size: 14px; font-weight: 500; white-space: nowrap; width: auto; }

.gb_Zd .gb_1d { -webkit-box-align: center; align-items: center; display: inline-flex; }

.gb_Zd .gb_r { fill: rgb(11, 87, 208); margin-left: 8px; }

.gb_Zd .gb_r circle { fill: rgb(255, 255, 255); }

.gb_Zd .gb_od .gb_Md { -webkit-box-flex: 1; flex-grow: 1; text-align: center; }

.gb_Zd .gb_od:hover { background: rgb(55, 99, 205); }

.gb_Zd .gb_od:hover .gb_r { fill: rgb(55, 99, 205); }

.gb_Zd .gb_od:focus, .gb_Zd .gb_od:active, .gb_Zd .gb_od:focus:hover { background: rgb(65, 106, 207); }

.gb_Zd .gb_od:focus .gb_r, .gb_Zd .gb_od:active .gb_r, .gb_Zd .gb_od:focus:hover .gb_r { fill: rgb(65, 106, 207); }

.gb_Zd .gb_od:hover, .gb_Zd .gb_od:focus, .gb_Zd .gb_od:active { box-shadow: rgba(66, 64, 67, 0.15) 0px 1px 3px 1px, rgba(60, 64, 67, 0.3) 0px 1px 2px 0px; }

.gb_Zd .gb_od:focus-visible { outline: rgb(65, 106, 207) solid 1px; outline-offset: 2px; }

.gb_Zd .gb_i.gb_od { background: rgb(168, 199, 250); color: rgb(6, 46, 111); }

.gb_Zd .gb_i.gb_od .gb_r { fill: rgb(168, 199, 250); }

.gb_Zd .gb_i.gb_od .gb_r circle { fill: rgb(6, 46, 111); }

.gb_Zd .gb_i.gb_od:hover { background: rgb(180, 203, 246); }

.gb_Zd .gb_i.gb_od:hover .gb_r { fill: rgb(180, 203, 246); }

.gb_Zd .gb_i.gb_od:focus, .gb_Zd .gb_i.gb_od:focus:hover, .gb_Zd .gb_i.gb_od:active { background: rgb(184, 205, 247); }

.gb_Zd .gb_i.gb_od:focus .gb_r, .gb_Zd .gb_i.gb_od:focus:hover .gb_r, .gb_Zd .gb_i.gb_od:active .gb_r { fill: rgb(184, 205, 247); }

.gb_Zd .gb_i.gb_od:focus-visible { outline-color: rgb(184, 205, 247); }

.gb_Zd .gb_i.gb_od:hover, .gb_Zd .gb_i.gb_od:focus, .gb_Zd .gb_i.gb_od:active { box-shadow: rgba(66, 64, 67, 0.15) 0px 1px 3px 1px, rgba(60, 64, 67, 0.3) 0px 1px 2px 0px; }

.gb_8c .gb_Xd, .gb_f .gb_Xd { float: right; }

.gb_d { padding: 8px; cursor: pointer; }

.gb_Pa .gb_oe:not(.gb_ka):focus img { background-color: rgba(0, 0, 0, 0.2); outline: none; border-radius: 50%; }

.gb_2d button svg, .gb_d { border-radius: 50%; }

.gb_2d button:focus:not(:focus-visible) svg, .gb_2d button:hover svg, .gb_2d button:active svg, .gb_d:focus:not(:focus-visible), .gb_d:hover, .gb_d:active, .gb_d[aria-expanded="true"] { outline: none; }

.gb_Rc .gb_2d.gb_xe button:focus-visible svg, .gb_2d button:focus-visible svg, .gb_d:focus-visible { outline: rgb(32, 33, 36) solid 1px; }

.gb_Rc .gb_2d button:focus-visible svg, .gb_Rc .gb_d:focus-visible { outline: rgb(241, 243, 244) solid 1px; }

@media (forced-colors: active) {
  .gb_Rc .gb_2d.gb_xe button:focus-visible svg, .gb_2d button:focus-visible svg, .gb_Rc .gb_2d button:focus-visible svg { outline: currentcolor solid 1px; }
}

.gb_Rc .gb_2d.gb_xe button:focus svg, .gb_Rc .gb_2d.gb_xe button:focus:hover svg, .gb_2d button:focus svg, .gb_2d button:focus:hover svg, .gb_d:focus, .gb_d:focus:hover { background-color: rgba(60, 64, 67, 0.1); }

.gb_Rc .gb_2d.gb_xe button:active svg, .gb_2d button:active svg, .gb_d:active { background-color: rgba(60, 64, 67, 0.12); }

.gb_Rc .gb_2d.gb_xe button:hover svg, .gb_2d button:hover svg, .gb_d:hover { background-color: rgba(60, 64, 67, 0.08); }

.gb_Da .gb_d.gb_Fa:hover { background-color: transparent; }

.gb_d[aria-expanded="true"], .gb_d:hover[aria-expanded="true"] { background-color: rgba(95, 99, 104, 0.24); }

.gb_d[aria-expanded="true"] .gb_h, .gb_d[aria-expanded="true"] .gb_5e { fill: rgb(95, 99, 104); opacity: 1; }

.gb_Rc .gb_2d button:hover svg, .gb_Rc .gb_d:hover { background-color: rgba(232, 234, 237, 0.08); }

.gb_Rc .gb_2d button:focus svg, .gb_Rc .gb_2d button:focus:hover svg, .gb_Rc .gb_d:focus, .gb_Rc .gb_d:focus:hover { background-color: rgba(232, 234, 237, 0.1); }

.gb_Rc .gb_2d button:active svg, .gb_Rc .gb_d:active { background-color: rgba(232, 234, 237, 0.12); }

.gb_Rc .gb_d[aria-expanded="true"], .gb_Rc .gb_d:hover[aria-expanded="true"] { background-color: rgba(255, 255, 255, 0.12); }

.gb_Rc .gb_d[aria-expanded="true"] .gb_h, .gb_Rc .gb_d[aria-expanded="true"] .gb_5e { fill: rgb(255, 255, 255); opacity: 1; }

.gb_Rd { padding: 4px; }

.gb_Pa.gb_Wd .gb_Rd { padding: 4px 2px; }

.gb_Pa.gb_Wd .gb_b.gb_Rd { padding-left: 6px; }

.gb_U { z-index: 991; line-height: normal; }

.gb_U.gb_3d { left: 0px; right: auto; }

@media (max-width: 350px) {
  .gb_U.gb_3d { left: 0px; }
}

.gb_4d .gb_U { top: 56px; }

.gb_S .gb_d, .gb_T .gb_S .gb_d { background-position: -64px -29px; }

.gb_y .gb_S .gb_d { background-position: -29px -29px; opacity: 1; }

.gb_S .gb_d, .gb_S .gb_d:hover, .gb_S .gb_d:focus { opacity: 1; }

.gb_md { display: none; }

@media screen and (max-width: 319px) {
  .gb_td:not(.gb_yd) .gb_S { display: none; visibility: hidden; }
}

.gb_l { display: none; }

.gb_gd { font-family: "Google Sans", Roboto, Helvetica, Arial, sans-serif; font-size: 20px; font-weight: 400; letter-spacing: 0.25px; line-height: 48px; margin-bottom: 2px; opacity: 1; overflow: hidden; padding-left: 16px; position: relative; text-overflow: ellipsis; vertical-align: middle; top: 2px; white-space: nowrap; -webkit-box-flex: 1; flex: 1 1 auto; }

.gb_gd.gb_hd { color: rgb(60, 64, 67); }

.gb_Pa.gb_Qa .gb_gd { margin-bottom: 0px; }

.gb_id.gb_jd .gb_gd { padding-left: 4px; }

.gb_Pa.gb_Qa .gb_kd { position: relative; top: -2px; }

.gb_Pa { color: black; min-width: 160px; position: relative; transition: box-shadow 250ms ease 0s; }

.gb_Pa.gb_0c { min-width: 120px; }

.gb_Pa.gb_rd .gb_sd { display: none; }

.gb_Pa.gb_rd .gb_td { height: 56px; }

header.gb_Pa { display: block; }

.gb_Pa svg { fill: currentcolor; }

.gb_ud { position: fixed; top: 0px; width: 100%; }

.gb_vd { box-shadow: rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px, rgba(0, 0, 0, 0.2) 0px 2px 4px -1px; }

.gb_wd { height: 64px; }

.gb_td { box-sizing: border-box; position: relative; width: 100%; display: flex; justify-content: space-between; min-width: min-content; }

.gb_Pa:not(.gb_Qa) .gb_td { padding: 8px; }

.gb_Pa.gb_xd .gb_td { -webkit-box-flex: 1; flex: 1 0 auto; }

.gb_Pa .gb_td.gb_yd.gb_zd { min-width: 0px; }

.gb_Pa.gb_Qa .gb_td { padding: 4px 4px 4px 8px; min-width: 0px; }

.gb_sd { height: 48px; vertical-align: middle; white-space: nowrap; -webkit-box-align: center; align-items: center; display: flex; user-select: none; }

.gb_Bd > .gb_sd { display: table-cell; width: 100%; }

.gb_id { padding-right: 30px; box-sizing: border-box; -webkit-box-flex: 1; flex: 1 0 auto; }

.gb_Pa.gb_Qa .gb_id { padding-right: 14px; }

.gb_Cd { -webkit-box-flex: 1; flex: 1 1 100%; }

.gb_Cd > :only-child { display: inline-block; }

.gb_Dd.gb_9c { padding-left: 4px; }

.gb_Dd.gb_Ed, .gb_Pa.gb_xd .gb_Dd, .gb_Pa.gb_Qa:not(.gb_f) .gb_Dd { padding-left: 0px; }

.gb_Pa.gb_Qa .gb_Dd.gb_Ed { padding-right: 0px; }

.gb_Pa.gb_Qa .gb_Dd.gb_Ed .gb_Da { margin-left: 10px; }

.gb_9c { display: inline; }

.gb_Pa.gb_3c .gb_Dd.gb_Fd, .gb_Pa.gb_f .gb_Dd.gb_Fd { padding-left: 2px; }

.gb_gd { display: inline-block; }

.gb_Dd { box-sizing: border-box; height: 48px; line-height: normal; padding: 0px 4px 0px 30px; -webkit-box-flex: 0; flex: 0 0 auto; justify-content: flex-end; }

.gb_f { height: 48px; }

.gb_Pa.gb_f { min-width: auto; }

.gb_f .gb_Dd { float: right; padding-left: 32px; }

.gb_f .gb_Dd.gb_Hd { padding-left: 0px; }

.gb_Id { font-size: 14px; max-width: 200px; overflow: hidden; padding: 0px 12px; text-overflow: ellipsis; white-space: nowrap; user-select: text; }

.gb_nd { transition: background-color 0.4s ease 0s; }

.gb_Nd { color: black; }

.gb_Rc { color: white; }

.gb_Pa a, .gb_Wc a { color: inherit; }

.gb_J { color: rgba(0, 0, 0, 0.87); }

.gb_Pa svg, .gb_Wc svg, .gb_id .gb_qd, .gb_8c .gb_qd { color: rgb(95, 99, 104); opacity: 1; }

.gb_Rc svg, .gb_Wc.gb_1c svg, .gb_Rc .gb_id .gb_qd, .gb_Rc .gb_id .gb_Qc, .gb_Rc .gb_id .gb_kd, .gb_Wc.gb_1c .gb_qd { color: rgba(255, 255, 255, 0.87); }

.gb_Rc .gb_id .gb_Pc:not(.gb_Od) { opacity: 0.87; }

.gb_hd { color: inherit; opacity: 1; text-rendering: optimizelegibility; -webkit-font-smoothing: antialiased; }

.gb_Rc .gb_hd, .gb_Nd .gb_hd { opacity: 1; }

.gb_Jd { position: relative; }

.gb_Kd { font-family: arial, sans-serif; line-height: normal; padding-right: 15px; }

a.gb_v, span.gb_v { color: rgba(0, 0, 0, 0.87); text-decoration: none; }

.gb_Rc a.gb_v, .gb_Rc span.gb_v { color: white; }

a.gb_v:focus { outline-offset: 2px; }

a.gb_v:hover { text-decoration: underline; }

.gb_w { display: inline-block; padding-left: 15px; }

.gb_w .gb_v { display: inline-block; line-height: 24px; vertical-align: middle; }

.gb_Pd { font-family: "Google Sans", Roboto, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; margin-left: 10px; margin-right: 8px; min-width: 96px; padding: 9px 23px; text-align: center; vertical-align: middle; border-radius: 4px; box-sizing: border-box; }

.gb_Pa.gb_f .gb_Pd { margin-left: 8px; }

#gb a.gb_oa.gb_Pd { cursor: pointer; }

.gb_oa.gb_Pd:hover { background: rgb(27, 102, 201); box-shadow: rgba(66, 64, 67, 0.15) 0px 1px 3px 1px, rgba(60, 64, 67, 0.3) 0px 1px 2px 0px; }

.gb_oa.gb_Pd:focus, .gb_oa.gb_Pd:hover:focus { background: rgb(28, 95, 186); box-shadow: rgba(66, 64, 67, 0.15) 0px 1px 3px 1px, rgba(60, 64, 67, 0.3) 0px 1px 2px 0px; }

.gb_oa.gb_Pd:active { background: rgb(27, 99, 193); box-shadow: rgba(66, 64, 67, 0.15) 0px 1px 3px 1px, rgba(60, 64, 67, 0.3) 0px 1px 2px 0px; }

.gb_Pd { background: rgb(26, 115, 232); border: 1px solid transparent; }

.gb_Pa.gb_Qa .gb_Pd { padding: 9px 15px; min-width: 80px; }

.gb_Ld { text-align: left; }

#gb .gb_Rc a.gb_Pd:not(.gb_i), #gb.gb_Rc a.gb_Pd:not(.gb_q) { background: rgb(255, 255, 255); border-color: rgb(218, 220, 224); box-shadow: none; color: rgb(26, 115, 232); }

#gb a.gb_oa.gb_i.gb_Pd { background: rgb(138, 180, 248); border: 1px solid transparent; box-shadow: none; color: rgb(32, 33, 36); }

#gb .gb_Rc a.gb_Pd:hover:not(.gb_i), #gb.gb_Rc a.gb_Pd:not(.gb_q):hover { background: rgb(248, 251, 255); border-color: rgb(204, 224, 252); }

#gb a.gb_oa.gb_i.gb_Pd:hover { background: rgb(147, 186, 249); border-color: transparent; box-shadow: rgba(0, 0, 0, 0.15) 0px 1px 3px 1px, rgba(0, 0, 0, 0.3) 0px 1px 2px; }

#gb .gb_Rc a.gb_Pd:focus:not(.gb_i), #gb .gb_Rc a.gb_Pd:focus:hover:not(.gb_i), #gb.gb_Rc a.gb_Pd:focus:not(.gb_i), #gb.gb_Rc a.gb_Pd:focus:hover:not(.gb_i) { background: rgb(244, 248, 255); outline: rgb(201, 221, 252) solid 1px; }

#gb a.gb_oa.gb_i.gb_Pd:focus, #gb a.gb_oa.gb_i.gb_Pd:focus:hover { background: rgb(166, 198, 250); border-color: transparent; box-shadow: none; }

#gb .gb_Rc a.gb_Pd:active:not(.gb_i), #gb.gb_Rc a.gb_Pd:not(.gb_q):active { background: rgb(236, 243, 254); }

#gb a.gb_oa.gb_i.gb_Pd:active { background: rgb(161, 195, 249); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.gb_Qd { display: none; }

@media screen and (max-width: 319px) {
  .gb_td:not(.gb_yd) .gb_S { display: none; visibility: hidden; }
}

.gb_Da { background-color: rgba(255, 255, 255, 0.88); border: 1px solid rgb(218, 220, 224); box-sizing: border-box; cursor: pointer; display: inline-block; max-height: 48px; overflow: hidden; outline: none; padding: 0px; vertical-align: middle; width: 134px; border-radius: 8px; }

.gb_Da.gb_i { background-color: transparent; border: 1px solid rgb(95, 99, 104); }

.gb_Ka { display: inherit; }

.gb_Da.gb_i .gb_Ka { background: rgb(255, 255, 255); border-radius: 4px; display: inline-block; left: 8px; margin-right: 5px; position: relative; padding: 3px; top: -1px; }

.gb_Da:hover { border: 1px solid rgb(210, 227, 252); background-color: rgba(248, 250, 255, 0.88); }

.gb_Da.gb_i:hover { background-color: rgba(241, 243, 244, 0.04); border: 1px solid rgb(95, 99, 104); }

.gb_Da:focus-visible, .gb_Da:focus { background-color: rgb(255, 255, 255); outline: rgb(32, 33, 36) solid 1px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.gb_Da.gb_i:focus-visible, .gb_Da.gb_i:focus { background-color: rgba(241, 243, 244, 0.12); outline: rgb(241, 243, 244) solid 1px; box-shadow: rgba(0, 0, 0, 0.15) 0px 1px 3px 1px, rgba(0, 0, 0, 0.3) 0px 1px 2px 0px; }

.gb_Da.gb_i:active, .gb_Da.gb_La.gb_i:focus { background-color: rgba(241, 243, 244, 0.1); border: 1px solid rgb(95, 99, 104); }

.gb_Ma { display: inline-block; padding-bottom: 2px; padding-left: 7px; padding-top: 2px; text-align: center; vertical-align: middle; line-height: 32px; width: 78px; }

.gb_Da.gb_i .gb_Ma { line-height: 26px; margin-left: 0px; padding-bottom: 0px; padding-left: 0px; padding-top: 0px; width: 72px; }

.gb_Ma.gb_Na { background-color: rgb(241, 243, 244); border-radius: 4px; margin-left: 8px; padding-left: 0px; line-height: 30px; }

.gb_Ma.gb_Na .gb_Oa { vertical-align: middle; }

.gb_Pa:not(.gb_Qa) .gb_Da { margin-left: 10px; margin-right: 4px; }

.gb_Ra { max-height: 32px; width: 78px; }

.gb_Da.gb_i .gb_Ra { max-height: 26px; width: 72px; }

.gb_k { background-size: 32px 32px; border: 0px; border-radius: 50%; display: block; margin: 0px; position: relative; height: 32px; width: 32px; z-index: 0; }

.gb_2a { background-color: rgb(232, 240, 254); border: 1px solid rgba(32, 33, 36, 0.08); position: relative; }

.gb_2a.gb_k { height: 30px; width: 30px; }

.gb_2a.gb_k:hover, .gb_2a.gb_k:active { box-shadow: none; }

.gb_3a { background: rgb(255, 255, 255); border: none; border-radius: 50%; bottom: 2px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; height: 14px; margin: 2px; position: absolute; right: 0px; width: 14px; }

.gb_4a { color: rgb(31, 113, 231); font: 400 22px / 32px "Google Sans", Roboto, Helvetica, Arial, sans-serif; text-align: center; text-transform: uppercase; }

@media (-webkit-min-device-pixel-ratio: 1.25), (min-resolution: 1.25dppx), (min-device-pixel-ratio:1.25) {
  .gb_k::before, .gb_5a::before { display: inline-block; transform: scale(0.5); transform-origin: left 0px; }
  .gb_A .gb_5a::before { }
}

.gb_k:hover, .gb_k:focus { box-shadow: rgba(0, 0, 0, 0.15) 0px 1px 0px; }

.gb_k:active { box-shadow: rgba(0, 0, 0, 0.15) 0px 2px 0px inset; }

.gb_k:active::after { background: rgba(0, 0, 0, 0.1); border-radius: 50%; content: ""; display: block; height: 100%; }

.gb_6a { cursor: pointer; line-height: 40px; min-width: 30px; opacity: 0.75; overflow: hidden; vertical-align: middle; text-overflow: ellipsis; }

.gb_d.gb_6a { width: auto; }

.gb_6a:hover, .gb_6a:focus { opacity: 0.85; }

.gb_7a .gb_6a, .gb_7a .gb_8a { line-height: 26px; }

#gb#gb.gb_7a a.gb_6a, .gb_7a .gb_8a { font-size: 11px; height: auto; }

.gb_9a { border-top: 4px solid rgb(0, 0, 0); border-left: 4px dashed transparent; border-right: 4px dashed transparent; display: inline-block; margin-left: 6px; opacity: 0.75; vertical-align: middle; }

.gb_Fa:hover .gb_9a { opacity: 0.85; }

.gb_Da > .gb_b { padding: 3px 3px 3px 4px; }

.gb_ab.gb_1a { color: rgb(255, 255, 255); }

.gb_y .gb_6a, .gb_y .gb_9a { opacity: 1; }

#gb#gb.gb_y.gb_y a.gb_6a, #gb#gb .gb_y.gb_y a.gb_6a { color: rgb(255, 255, 255); }

.gb_y.gb_y .gb_9a { border-top-color: rgb(255, 255, 255); opacity: 1; }

.gb_T .gb_k:hover, .gb_y .gb_k:hover, .gb_T .gb_k:focus, .gb_y .gb_k:focus { box-shadow: rgba(0, 0, 0, 0.15) 0px 1px 0px, rgba(0, 0, 0, 0.2) 0px 1px 2px; }

.gb_bb .gb_b, .gb_cb .gb_b { position: absolute; right: 1px; }

.gb_b.gb_x, .gb_db.gb_x, .gb_Fa.gb_x { -webkit-box-flex: 0; flex: 0 1 auto; }

.gb_eb.gb_fb .gb_6a { width: 30px !important; }

.gb_j { height: 40px; position: absolute; right: -5px; top: -5px; width: 40px; }

.gb_gb .gb_j, .gb_hb .gb_j { right: 0px; top: 0px; }

.gb_b .gb_d { padding: 4px; }

.gb_n { display: none; }

sentinel { }
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/css
Content-Transfer-Encoding: binary
Content-Location: https://fonts.googleapis.com/css?family=Google+Sans_old:300,400,500,700

@charset "utf-8";

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiIUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+308, U+530-58F, U+2010, U+2024, U+25CC, U+FB13-FB17; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjMUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+900-97F, U+1CD0-1CF9, U+200C-200D, U+20A8, U+20B9, U+25CC, U+A830-A839, U+A8E0-A8FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPi0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+589, U+10A0-10FF, U+1C90-1CBA, U+1CBD-1CBF, U+2D00-2D2F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPhEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+A01-A76, U+200C-200D, U+20B9, U+25CC, U+262C, U+A830-A839; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjAUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+590-5FF, U+200C-2010, U+20AA, U+25CC, U+FB1D-FB4F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjsUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E81-EDF, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiQUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+B82-BFA, U+200C-200D, U+20B9, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E01-E5B, U+200C-200D, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPj0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjwUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 400; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjIUvbQoi-E.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiIUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+308, U+530-58F, U+2010, U+2024, U+25CC, U+FB13-FB17; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjMUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+900-97F, U+1CD0-1CF9, U+200C-200D, U+20A8, U+20B9, U+25CC, U+A830-A839, U+A8E0-A8FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPi0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+589, U+10A0-10FF, U+1C90-1CBA, U+1CBD-1CBF, U+2D00-2D2F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPhEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+A01-A76, U+200C-200D, U+20B9, U+25CC, U+262C, U+A830-A839; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjAUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+590-5FF, U+200C-2010, U+20AA, U+25CC, U+FB1D-FB4F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjsUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E81-EDF, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiQUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+B82-BFA, U+200C-200D, U+20B9, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E01-E5B, U+200C-200D, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPj0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjwUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 500; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjIUvbQoi-E.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiIUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+308, U+530-58F, U+2010, U+2024, U+25CC, U+FB13-FB17; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+301, U+400-45F, U+490-491, U+4B0-4B1, U+2116; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjMUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+900-97F, U+1CD0-1CF9, U+200C-200D, U+20A8, U+20B9, U+25CC, U+A830-A839, U+A8E0-A8FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPi0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+589, U+10A0-10FF, U+1C90-1CBA, U+1CBD-1CBF, U+2D00-2D2F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+370-3FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPhEUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+A01-A76, U+200C-200D, U+20B9, U+25CC, U+262C, U+A830-A839; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjAUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+590-5FF, U+200C-2010, U+20AA, U+25CC, U+FB1D-FB4F; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjsUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E81-EDF, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiQUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+964-965, U+B82-BFA, U+200C-200D, U+20B9, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPiYUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+E01-E5B, U+200C-200D, U+25CC; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPj0UvbQoi-Entw.woff2") format("woff2"); unicode-range: U+102-103, U+110-111, U+128-129, U+168-169, U+1A0-1A1, U+1AF-1B0, U+300-301, U+303-304, U+308-309, U+323, U+329, U+1EA0-1EF9, U+20AB; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjwUvbQoi-Entw.woff2") format("woff2"); unicode-range: U+100-2AF, U+304, U+308, U+329, U+1E00-1E9F, U+1EF2-1EFF, U+2020, U+20A0-20AB, U+20AD-20CF, U+2113, U+2C60-2C7F, U+A720-A7FF; }

@font-face { font-family: "Google Sans"; font-style: normal; font-weight: 700; src: url("https://fonts.gstatic.com/s/googlesans/v46/4UasrENHsxJlGDuGo1OIlJfC6l_24rlCK1Yo_Iqcsih3SAyH6cAwhX9RPjIUvbQoi-E.woff2") format("woff2"); unicode-range: U+0-FF, U+131, U+152-153, U+2BB-2BC, U+2C6, U+2DA, U+2DC, U+304, U+308, U+329, U+2000-206F, U+2074, U+20AC, U+2122, U+2191, U+2193, U+2212, U+2215, U+FEFF, U+FFFD; }
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/css
Content-Transfer-Encoding: binary
Content-Location: https://www.gstatic.com/_/apps-fileview/_/ss/k=apps-fileview.v.omJv0zZNxLk.L.W.O/am=AAAE/d=0/rs=AO0039tfU3F6Yks5o2y0ftEU4qi8duRDBA

@charset "utf-8";

@keyframes shimmer { 
  0% { background-position: 100% 50%; }
  100% { background-position: 0px 50%; }
}

@keyframes fadeInAnimation { 
  0% { opacity: 0; }
  100% { opacity: 1; }
}

.ja0jmf { align-content: center; animation: 200ms ease 0s 1 normal none running fadeInAnimation; background-color: var(--dt-surface,#fff); display: flex; flex-direction: column; height: 100%; position: absolute; top: 0px; width: 100%; z-index: 3000; }

.F6wkof { animation: 2.2s ease 0s infinite normal none running shimmer; background-image: ; background-position-x: ; background-position-y: ; background-size: ; background-repeat-x: ; background-repeat-y: ; background-attachment: ; background-origin: ; background-clip: ; background-color: var(--dt-inverse-on-surface,#dadce0); }

@media (forced-colors: active) {
  .F6wkof { border: 1px solid var(--dt-outline,#80868b); }
}

.HrDxdd { border-radius: 1rem; height: 1rem; margin-left: 1rem; margin-top: 0.5rem; }

.HrDxdd:nth-child(2n+1) { margin-top: 1.5rem; }

.ISv2N { background-color: transparent; border: none; color: inherit; cursor: pointer; fill: currentcolor; margin-right: 1rem; margin-top: 0.125rem; outline: none; padding: 0.75rem; text-decoration: none; }

.EebkFb { align-items: center; border-bottom: 1px solid var(--dt-outline,#80868b); display: flex; justify-content: space-between; margin-bottom: 1rem; margin-top: 0.3125rem; padding-bottom: 0.375rem; width: 100%; }

.gAm2E { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); color: var(--dt-on-background,#3c4043); margin-left: 20px; }

.NFRm8d { align-items: center; animation: 200ms ease 0s 1 normal none running fadeInAnimation; background-color: var(--dt-surface,#fff); display: flex; flex-direction: column; height: 100%; width: 100%; z-index: 3000; }

.C4MDDc { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,0.025em); color: var(--dt-on-surface,#3c4043); margin-top: 5.125rem; }

.Q6yead { fill: currentcolor; overflow: hidden; }

.mig17c { overflow: visible; }

[dir="rtl"] .Q6yead.wSyMnf { transform: scaleX(-1); }

@media (forced-colors: active) {
  .Q6yead.QJZfhe.QJZfhe { fill: canvastext; }
}

.A5Gtre { font-style: inherit; font-variant: inherit; font-stretch: inherit; line-height: inherit; font-family: inherit; font-optical-sizing: inherit; font-kerning: inherit; font-feature-settings: inherit; font-variation-settings: inherit; font-size: 100%; font-weight: inherit; text-decoration: none; }

.A5Gtre:hover, .A5Gtre:active, .A5Gtre:focus { text-decoration: underline; }

.cS0c5e { clip-path: inset(50%); clip: rect(1px, 1px, 1px, 1px); height: 1px; margin: -1px; opacity: 0; overflow: hidden; padding: 0px; position: absolute; width: 1px; }

.VIpgJd-TzA9Ye-eEGnhe { position: relative; display: inline-block; }

* html .VIpgJd-TzA9Ye-eEGnhe { display: inline; }

:first-child + html .VIpgJd-TzA9Ye-eEGnhe { display: inline; }

.tk3N6e-VCkuzd { box-shadow: rgba(0, 0, 0, 0.2) 0px 1px 3px; background-color: rgb(255, 255, 255); border-width: 1px; border-style: solid; border-image: initial; border-color: rgb(187, 187, 187) rgb(187, 187, 187) rgb(168, 168, 168); padding: 16px; position: absolute; z-index: 1201 !important; }

.tk3N6e-VCkuzd-kmh2Gb { background: url("//ssl.gstatic.com/ui/v1/icons/common/x_8px.png") no-repeat; border: 1px solid transparent; height: 21px; opacity: 0.4; outline: 0px; position: absolute; right: 2px; top: 2px; width: 21px; }

.tk3N6e-VCkuzd-kmh2Gb:focus { border: 1px solid rgb(77, 144, 254); opacity: 0.8; }

.tk3N6e-VCkuzd-hFsbo { position: absolute; }

.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc, .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { display: block; height: 0px; position: absolute; width: 0px; }

.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc { border: 9px solid; }

.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border: 8px solid; }

.tk3N6e-VCkuzd-Ya1KTb { bottom: 0px; }

.tk3N6e-VCkuzd-d6mlqf { top: -9px; }

.tk3N6e-VCkuzd-y6n2Me { left: -9px; }

.tk3N6e-VCkuzd-cX0Lwc { right: 0px; }

.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc, .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { left: -9px; }

.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc { border-bottom-width: 0px; }

.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG, .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG { border-color: rgb(255, 255, 255) transparent; left: -8px; }

.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG { border-bottom-width: 0px; }

.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { border-top-width: 0px; }

.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG { border-top-width: 0px; top: 1px; }

.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc, .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc { border-color: transparent rgb(187, 187, 187); top: -9px; }

.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG, .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG { border-color: transparent rgb(255, 255, 255); top: -8px; }

.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc { border-left-width: 0px; }

.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG { border-left-width: 0px; left: 1px; }

.tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc, .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG { border-right-width: 0px; }

.tk3N6e-suEOdc { border-radius: 0px; box-shadow: none; background-color: rgb(42, 42, 42); border: 1px solid rgb(255, 255, 255); color: rgb(255, 255, 255); cursor: default; display: block; margin-left: -1px; opacity: 1; padding: 7px 9px; position: absolute; visibility: visible; white-space: pre-wrap; word-break: break-word; }

.tk3N6e-suEOdc-ZYIfFd { opacity: 0; visibility: hidden; left: 20px !important; top: 20px !important; }

.tk3N6e-suEOdc-wZVHld { display: none; }

.tk3N6e-suEOdc-hFsbo { pointer-events: none; position: absolute; }

.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { content: ""; display: block; height: 0px; position: absolute; width: 0px; }

.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc { border: 6px solid; }

.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { border: 5px solid; }

.tk3N6e-suEOdc-Ya1KTb { bottom: 0px; }

.tk3N6e-suEOdc-d6mlqf { top: -6px; }

.tk3N6e-suEOdc-y6n2Me { left: -6px; }

.tk3N6e-suEOdc-cX0Lwc { right: 0px; }

.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc { border-color: rgb(255, 255, 255) transparent; left: -6px; }

.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG, .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-color: rgb(42, 42, 42) transparent; left: -5px; }

.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG { border-bottom-width: 0px; }

.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc { border-top-width: 0px; }

.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-top-width: 0px; top: 1px; }

.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc { border-color: transparent rgb(255, 255, 255); top: -6px; }

.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG, .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG { border-color: transparent rgb(42, 42, 42); top: -5px; }

.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc { border-left-width: 0px; }

.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG { border-left-width: 0px; left: 1px; }

.tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG { border-right-width: 0px; }

.cAHxfe { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); background: var(--dt-inverse-surface,rgb(32,33,36)); border-radius: 0.25rem; border: 1px solid transparent; box-sizing: border-box; color: var(--dt-inverse-on-surface,rgb(218,220,224)); margin: 0px; max-width: 100vw; min-height: 1.375rem; min-width: 3.5rem; padding: 0.25rem 0.5rem; text-align: center; z-index: 6000; }

.cAHxfe:not(.tk3N6e-suEOdc-ZYIfFd) { opacity: 1; transform: scale(1); }

.cAHxfe.tk3N6e-suEOdc-ZYIfFd { opacity: 0; transform: scale(0.9); width: 0px; }

.cAHxfe .tk3N6e-suEOdc-hFsbo { display: none; }

.pDtC4e { display: inline-block; }

.yYWAMb { background: var(--dt-background,#fff); color: var(--dt-on-background,rgb(60,64,67)); }

.XV0XSd { --dt-display-1-font: 400 4rem/4.75rem "Google Sans Display"; --dt-display-1-spacing: 0; --dt-display-large-font: 400 3.5rem/4rem "Google Sans Display"; --dt-display-large-spacing: 0; --dt-display-medium-font: 400 2.75rem/3.25rem "Google Sans Display"; --dt-display-medium-spacing: 0; --dt-display-small-font: 400 2.25rem/2.75rem "Google Sans"; --dt-display-small-spacing: 0; --dt-headline-large-font: 400 2rem/2.5rem "Google Sans"; --dt-headline-large-spacing: 0; --dt-headline-medium-font: 400 1.75rem/2.25rem "Google Sans"; --dt-headline-medium-spacing: 0; --dt-headline-small-font: 400 1.5rem/2rem "Google Sans"; --dt-headline-small-spacing: 0; --dt-title-large-font: 400 1.375rem/1.75rem "Google Sans"; --dt-title-large-spacing: 0; --dt-headline-6-font: 400 1.125rem/1.5rem "Google Sans"; --dt-headline-6-spacing: 0; --dt-title-medium-font: 500 1rem/1.5rem "Google Sans"; --dt-title-medium-spacing: 0.00625em; --dt-title-small-font: 500 0.875rem/1.25rem "Google Sans"; --dt-title-small-spacing: 0.0178571429em; --dt-subtitle-1-font: 500 1rem/1.5rem "Roboto"; --dt-subtitle-1-spacing: 0.0125em; --dt-label-large-font: 500 0.875rem/1.25rem "Roboto"; --dt-label-large-spacing: 0.0178571429em; --dt-label-medium-font: 500 0.75rem/1rem "Roboto"; --dt-label-medium-spacing: 0.0208333333em; --dt-label-small-font: 500 0.6875rem/1rem "Roboto"; --dt-label-small-spacing: 0.0727272727em; --dt-label-small-transform: uppercase; --dt-body-large-font: 400 1rem/1.5rem "Roboto"; --dt-body-large-spacing: 0.00625em; --dt-body-medium-font: 400 0.875rem/1.25rem "Roboto"; --dt-body-medium-spacing: 0.0142857143em; --dt-body-small-font: 400 0.75rem/1rem "Roboto"; --dt-body-small-spacing: 0.025em; --dt-corner-banner: 0.25rem; --dt-corner-button: 0.25rem; --dt-corner-card: 0.375rem; --dt-corner-card-thumbnail: 0; --dt-corner-chip: 6.25rem; --dt-corner-chip-avatar: 6.25rem; --dt-corner-chip-suggestive: 0.5rem; --dt-corner-dialog: 0.5rem; --dt-corner-dialog-anchored: 0.5rem; --dt-corner-fab: 6.25rem; --dt-corner-fab-large: 6.25rem; --dt-corner-field: 0.375rem; --dt-corner-field-filled: 0.375rem 0.375rem 0 0; --dt-corner-field-search: 0.5rem; --dt-corner-icon-button: 6.25rem; --dt-corner-landmark: 0; --dt-corner-menu: 0.25rem; --dt-corner-mole: 0.25rem; --dt-corner-nav-drawer: 0 1.5rem 1.5rem 0; --dt-corner-region: 0.5rem; --dt-corner-tile: 0.375rem; }

.vhoiae, .X9XeLb, .cWKK1c, .aJfoSc, .TOb6Ze { --dt-display-1-font: 400 3.5625rem/4rem "Google Sans"; --dt-display-1-spacing: 0; --dt-display-large-font: 400 3.5625rem/4rem "Google Sans"; --dt-display-large-spacing: 0; --dt-display-medium-font: 400 2.8125rem/3.25rem "Google Sans"; --dt-display-medium-spacing: 0; --dt-display-small-font: 400 2.25rem/2.75rem "Google Sans"; --dt-display-small-spacing: 0; --dt-headline-large-font: 400 2rem/2.5rem "Google Sans"; --dt-headline-large-spacing: 0; --dt-headline-medium-font: 400 1.75rem/2.25rem "Google Sans"; --dt-headline-medium-spacing: 0; --dt-headline-small-font: 400 1.5rem/2rem "Google Sans"; --dt-headline-small-spacing: 0; --dt-title-large-font: 400 1.375rem/1.75rem "Google Sans"; --dt-title-large-spacing: 0; --dt-headline-6-font: 400 1.375rem/1.75rem "Google Sans"; --dt-headline-6-spacing: 0; --dt-title-medium-font: 500 1rem/1.5rem "Google Sans Text"; --dt-title-medium-spacing: 0; --dt-title-small-font: 500 0.875rem/1.25rem "Google Sans Text"; --dt-title-small-spacing: 0; --dt-subtitle-1-font: 500 1rem/1.5rem "Google Sans Text"; --dt-subtitle-1-spacing: 0; --dt-label-large-font: 500 0.875rem/1.25rem "Google Sans Text"; --dt-label-large-spacing: 0; --dt-label-medium-font: 500 0.75rem/1rem "Google Sans Text"; --dt-label-medium-spacing: 0; --dt-label-small-font: 500 0.6875rem/1rem "Google Sans Text"; --dt-label-small-spacing: 0.0090909091em; --dt-label-small-transform: none; --dt-body-large-font: 400 1rem/1.5rem "Google Sans Text"; --dt-body-large-spacing: 0; --dt-body-medium-font: 400 0.875rem/1.25rem "Google Sans Text"; --dt-body-medium-spacing: 0; --dt-body-small-font: 400 0.75rem/1rem "Google Sans Text"; --dt-body-small-spacing: 0.0083333333em; --dt-corner-banner: 0.5rem; --dt-corner-button: 6.25rem; --dt-corner-card: 0.75rem; --dt-corner-card-thumbnail: 0.25rem; --dt-corner-chip: 0.5rem; --dt-corner-chip-avatar: 6.25rem; --dt-corner-chip-suggestive: 0.5rem; --dt-corner-dialog: 0.5rem; --dt-corner-dialog-anchored: 0.5rem; --dt-corner-fab: 1rem; --dt-corner-fab-large: 1.75rem; --dt-corner-field: 0.25rem; --dt-corner-field-filled: 0.25rem 0.25rem 0 0; --dt-corner-field-search: 0.25rem; --dt-corner-icon-button: 6.25rem; --dt-corner-landmark: 1rem; --dt-corner-menu: 0.25rem; --dt-corner-mole: 1rem; --dt-corner-nav-drawer: 6.25rem; --dt-corner-region: 0.75rem; --dt-corner-tile: 1rem; }

.vhoiae .tk3N6e-suEOdc, .X9XeLb .tk3N6e-suEOdc, .cWKK1c .tk3N6e-suEOdc, .aJfoSc .tk3N6e-suEOdc, .TOb6Ze .tk3N6e-suEOdc { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); background: var(--dt-inverse-surface,rgb(32,33,36)); border-radius: 0.25rem; border: 1px solid transparent; box-sizing: border-box; color: var(--dt-inverse-on-surface,rgb(218,220,224)); margin: 0px; max-width: 100vw; min-height: 1.375rem; min-width: 3.5rem; padding: 0.25rem 0.5rem; text-align: center; z-index: 6000; }

.vhoiae .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd), .X9XeLb .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd), .cWKK1c .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd), .aJfoSc .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd), .TOb6Ze .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd) { opacity: 1; transform: scale(1); }

.vhoiae .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd, .X9XeLb .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd, .cWKK1c .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd, .aJfoSc .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd, .TOb6Ze .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd { opacity: 0; transform: scale(0.9); width: 0px; }

.vhoiae .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo, .X9XeLb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo, .cWKK1c .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo, .aJfoSc .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo, .TOb6Ze .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo { display: none; }

.vhoiae .XKSfm-Sx9Kwc, .X9XeLb .XKSfm-Sx9Kwc, .cWKK1c .XKSfm-Sx9Kwc, .aJfoSc .XKSfm-Sx9Kwc, .TOb6Ze .XKSfm-Sx9Kwc { background-color: var(--dt-surface,#fff); border-radius: var(--dt-corner-dialog,.5rem); color: var(--dt-on-surface,rgb(60,64,67)); }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); background-color: var(--dt-surface,#fff); }

.vhoiae .XKSfm-Sx9Kwc-r4nke, .X9XeLb .XKSfm-Sx9Kwc-r4nke, .cWKK1c .XKSfm-Sx9Kwc-r4nke, .aJfoSc .XKSfm-Sx9Kwc-r4nke, .TOb6Ze .XKSfm-Sx9Kwc-r4nke { background-color: var(--dt-surface,#fff); }

.vhoiae .XKSfm-Sx9Kwc-r4nke-TvD9Pc, .X9XeLb .XKSfm-Sx9Kwc-r4nke-TvD9Pc, .cWKK1c .XKSfm-Sx9Kwc-r4nke-TvD9Pc, .aJfoSc .XKSfm-Sx9Kwc-r4nke-TvD9Pc, .TOb6Ze .XKSfm-Sx9Kwc-r4nke-TvD9Pc { color: var(--dt-on-surface,rgb(60,64,67)); }

.vhoiae .XKSfm-Sx9Kwc-r4nke-fmcmS, .X9XeLb .XKSfm-Sx9Kwc-r4nke-fmcmS, .cWKK1c .XKSfm-Sx9Kwc-r4nke-fmcmS, .aJfoSc .XKSfm-Sx9Kwc-r4nke-fmcmS, .TOb6Ze .XKSfm-Sx9Kwc-r4nke-fmcmS { font: var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-headline-small-spacing,0); }

.vhoiae .XKSfm-Sx9Kwc-dI4VCc, .X9XeLb .XKSfm-Sx9Kwc-dI4VCc, .cWKK1c .XKSfm-Sx9Kwc-dI4VCc, .aJfoSc .XKSfm-Sx9Kwc-dI4VCc, .TOb6Ze .XKSfm-Sx9Kwc-dI4VCc { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); background-color: var(--dt-surface,#fff); border-color: var(--dt-outline,rgb(128,134,139)); border-radius: var(--dt-corner-field,.375rem); box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); height: 2.625rem; }

.vhoiae .XKSfm-Sx9Kwc-dI4VCc:focus, .X9XeLb .XKSfm-Sx9Kwc-dI4VCc:focus, .cWKK1c .XKSfm-Sx9Kwc-dI4VCc:focus, .aJfoSc .XKSfm-Sx9Kwc-dI4VCc:focus, .TOb6Ze .XKSfm-Sx9Kwc-dI4VCc:focus { border-color: var(--dt-primary,rgb(26,115,232)); border-width: 0.125rem; box-shadow: none; }

.vhoiae .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc, .X9XeLb .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc, .cWKK1c .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc, .aJfoSc .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc, .TOb6Ze .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { background: none; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,.0178571429em); overflow: visible; border-radius: var(--dt-corner-button,.25rem); color: var(--dt-primary,rgb(26,115,232)); text-transform: capitalize; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button::after, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after { transition: color 15ms linear 0s, background 15ms linear 0s, opacity 15ms linear 0s; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover { box-shadow: none; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before { background-color: currentcolor; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.12; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.08; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::after, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after { bottom: 0px; border-radius: 0.375rem; content: ""; display: block; height: 100%; left: 0px; outline: solid 2px var(--dt-primary,rgb(26,115,232)); outline-offset: 3px; position: absolute; width: 100%; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc { overflow: visible; background-color: var(--dt-primary,rgb(26,115,232)); color: var(--dt-on-primary,#fff); }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after { transition: color 15ms linear 0s, background 15ms linear 0s, opacity 15ms linear 0s; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover { box-shadow: none; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before { background-color: currentcolor; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.12; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.08; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after { bottom: 0px; border-radius: 0.375rem; content: ""; display: block; height: 100%; left: 0px; outline: solid 2px var(--dt-primary,rgb(26,115,232)); outline-offset: 3px; position: absolute; width: 100%; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe { padding-top: 0.3125rem; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc { background-color: var(--dt-surface,#fff); background-image: none; border: .0625rem solid var(--dt-outline,rgb(128,134,139)); box-shadow: none; box-sizing: border-box; color: var(--dt-primary,rgb(26,115,232)); }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover { border: .0625rem solid var(--dt-outline,rgb(128,134,139)); box-shadow: none; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me) { overflow: visible; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me), .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after { transition: color 15ms linear 0s, background 15ms linear 0s, opacity 15ms linear 0s; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover { box-shadow: none; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before { background-color: currentcolor; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.12; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before { border-radius: var(--dt-corner-button,.25rem); opacity: 0.08; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after { bottom: 0px; border-radius: 0.375rem; content: ""; display: block; height: 100%; left: 0px; outline: solid 2px var(--dt-primary,rgb(26,115,232)); outline-offset: 3px; position: absolute; width: 100%; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me { color: var(--dt-on-background,rgb(60,64,67)); opacity: 0.38; }

.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before, .TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before { background-color: inherit; }

.vhoiae ::-webkit-scrollbar, .X9XeLb ::-webkit-scrollbar, .cWKK1c ::-webkit-scrollbar, .aJfoSc ::-webkit-scrollbar, .TOb6Ze ::-webkit-scrollbar { height: 8px; width: 8px; }

.vhoiae ::-webkit-scrollbar-corner, .X9XeLb ::-webkit-scrollbar-corner, .cWKK1c ::-webkit-scrollbar-corner, .aJfoSc ::-webkit-scrollbar-corner, .TOb6Ze ::-webkit-scrollbar-corner { background: transparent; }

.vhoiae ::-webkit-scrollbar-thumb, .X9XeLb ::-webkit-scrollbar-thumb, .cWKK1c ::-webkit-scrollbar-thumb, .aJfoSc ::-webkit-scrollbar-thumb, .TOb6Ze ::-webkit-scrollbar-thumb { background-clip: padding-box; background-color: var(--dt-outline-variant,rgb(218,220,224)); border-radius: 100px; border: none; height: 8px; padding: 100px 0px 0px; width: 8px; }

.vhoiae ::-webkit-scrollbar-thumb:hover, .X9XeLb ::-webkit-scrollbar-thumb:hover, .cWKK1c ::-webkit-scrollbar-thumb:hover, .aJfoSc ::-webkit-scrollbar-thumb:hover, .TOb6Ze ::-webkit-scrollbar-thumb:hover { background-color: var(--dt-outline,rgb(128,134,139)); }

.vhoiae ::-webkit-scrollbar-thumb:active, .X9XeLb ::-webkit-scrollbar-thumb:active, .cWKK1c ::-webkit-scrollbar-thumb:active, .aJfoSc ::-webkit-scrollbar-thumb:active, .TOb6Ze ::-webkit-scrollbar-thumb:active { background-color: var(--dt-outline,rgb(128,134,139)); }

.vhoiae ::-webkit-scrollbar-track, .X9XeLb ::-webkit-scrollbar-track, .cWKK1c ::-webkit-scrollbar-track, .aJfoSc ::-webkit-scrollbar-track, .TOb6Ze ::-webkit-scrollbar-track { background-color: transparent; border: none; box-shadow: none; height: 8px; width: 8px; }

.vhoiae ::-webkit-scrollbar-track:hover, .X9XeLb ::-webkit-scrollbar-track:hover, .cWKK1c ::-webkit-scrollbar-track:hover, .aJfoSc ::-webkit-scrollbar-track:hover, .TOb6Ze ::-webkit-scrollbar-track:hover { border: none; box-shadow: none; }

@media (forced-colors: active) {
  .vhoiae ::-webkit-scrollbar-thumb, .vhoiae ::-webkit-scrollbar-thumb:hover, .vhoiae ::-webkit-scrollbar-thumb:active, .X9XeLb ::-webkit-scrollbar-thumb, .X9XeLb ::-webkit-scrollbar-thumb:hover, .X9XeLb ::-webkit-scrollbar-thumb:active, .cWKK1c ::-webkit-scrollbar-thumb, .cWKK1c ::-webkit-scrollbar-thumb:hover, .cWKK1c ::-webkit-scrollbar-thumb:active, .aJfoSc ::-webkit-scrollbar-thumb, .aJfoSc ::-webkit-scrollbar-thumb:hover, .aJfoSc ::-webkit-scrollbar-thumb:active, .TOb6Ze ::-webkit-scrollbar-thumb, .TOb6Ze ::-webkit-scrollbar-thumb:hover, .TOb6Ze ::-webkit-scrollbar-thumb:active { background-color: canvastext; }
}

.XV0XSd.KkxPLb { --dt-background: #fff; --dt-on-background: rgb(60,64,67); --dt-on-background-secondary: rgb(95,99,104); --dt-outline: rgb(128,134,139); --dt-outline-variant: rgb(218,220,224); --dt-on-disabled: rgba(60,64,67,0.38); --dt-disabled: rgba(60,64,67,0.12); --dt-inverse-on-surface: rgb(218,220,224); --dt-inverse-surface: rgb(32,33,36); --dt-on-surface-variant: rgb(95,99,104); --dt-on-surface-secondary: rgb(95,99,104); --dt-on-surface: rgb(60,64,67); --dt-surface-tint: rgb(241,243,244); --dt-surface-variant: rgb(241,243,244); --dt-surface1: #fff; --dt-surface1-shadow: 0 1px 2px 0 rgba(60,64,67,0.3),0 1px 3px 1px rgba(60,64,67,0.15); --dt-surface2: #fff; --dt-surface2-shadow: 0 1px 2px 0 rgba(60,64,67,0.3),0 2px 6px 2px rgba(60,64,67,0.15); --dt-surface3: #fff; --dt-surface3-shadow: 0 1px 3px 0 rgba(60,64,67,0.3),0 4px 8px 3px rgba(60,64,67,0.15); --dt-surface4: #fff; --dt-surface4-shadow: 0 2px 3px 0 rgba(60,64,67,0.3),0 6px 10px 4px rgba(60,64,67,0.15); --dt-surface5: #fff; --dt-surface5-shadow: 0 4px 4px 0 rgba(60,64,67,0.3),0 8px 12px 6px rgba(60,64,67,0.15); --dt-surface: #fff; --dt-scrim: rgba(32,33,36,0.6); --dt-scrim-2x: rgb(32,33,36); --dt-on-primary-container: rgb(60,64,67); --dt-on-primary: #fff; --dt-primary-action-state-layer: rgb(25,103,210); --dt-primary-action-stateful: rgb(24,90,188); --dt-primary-action: rgb(25,103,210); --dt-primary-container-icon: rgb(25,103,210); --dt-primary-container-link: rgb(25,103,210); --dt-primary-container: rgb(232,240,254); --dt-primary-icon: #fff; --dt-primary-link: #fff; --dt-primary-outline: rgb(24,90,188); --dt-primary: rgb(26,115,232); --dt-on-secondary-container: rgb(60,64,67); --dt-on-secondary: #fff; --dt-secondary-action-state-layer: rgb(60,64,67); --dt-secondary-action-stateful: rgb(32,33,36); --dt-secondary-action: rgb(60,64,67); --dt-secondary-container-icon: rgb(60,64,67); --dt-secondary-container-link: rgb(25,103,210); --dt-secondary-container: rgb(241,243,244); --dt-secondary-icon: #fff; --dt-secondary-link: #fff; --dt-secondary-outline: rgb(60,64,67); --dt-secondary: rgb(60,64,67); --dt-on-tertiary-container: rgb(60,64,67); --dt-on-tertiary: #fff; --dt-tertiary-action-state-layer: rgb(19,115,51); --dt-tertiary-action-stateful: rgb(13,101,45); --dt-tertiary-action: rgb(19,115,51); --dt-tertiary-container-icon: rgb(19,115,51); --dt-tertiary-container-link: rgb(19,115,51); --dt-tertiary-container: rgb(230,244,234); --dt-tertiary-icon: #fff; --dt-tertiary-link: #fff; --dt-tertiary-outline: rgb(19,115,51); --dt-tertiary: rgb(24,128,56); --dt-on-neutral-container: rgb(60,64,67); --dt-on-neutral: #fff; --dt-neutral-action-state-layer: rgb(60,64,67); --dt-neutral-action-stateful: rgb(32,33,36); --dt-neutral-action: rgb(60,64,67); --dt-neutral-container-icon: rgb(60,64,67); --dt-neutral-container-link: rgb(25,103,210); --dt-neutral-container: rgb(241,243,244); --dt-neutral-icon: #fff; --dt-neutral-link: #fff; --dt-neutral-outline: rgb(60,64,67); --dt-neutral: rgb(60,64,67); --dt-error-action-state-layer: rgb(197,34,31); --dt-error-action-stateful: rgb(179,20,18); --dt-error-action: rgb(197,34,31); --dt-error-container-icon: rgb(197,34,31); --dt-error-container-link: rgb(197,34,31); --dt-error-container: rgb(252,232,230); --dt-error-icon: #fff; --dt-error-link: #fff; --dt-error-outline: rgb(179,20,18); --dt-error: rgb(217,48,37); --dt-on-error-container: rgb(60,64,67); --dt-on-error: #fff; --dt-on-warning-container: rgb(60,64,67); --dt-on-warning: rgb(32,33,36); --dt-warning-action-state-layer: rgb(234,134,0); --dt-warning-action-stateful: rgb(32,33,36); --dt-warning-action: rgb(60,64,67); --dt-warning-container-icon: rgb(60,64,67); --dt-warning-container-link: rgb(60,64,67); --dt-warning-container: rgb(254,247,224); --dt-warning-icon: rgb(60,64,67); --dt-warning-link: rgb(60,64,67); --dt-warning-outline: rgb(234,134,0); --dt-warning: rgb(249,171,0); --gm3-sys-color-background: #fff; --gm3-sys-color-background-rgb: 255,255,255; --gm3-sys-color-error: #b3261e; --gm3-sys-color-error-rgb: 179,38,30; --gm3-sys-color-error-container: #f9dedc; --gm3-sys-color-error-container-rgb: 249,222,220; --gm3-sys-color-inverse-on-surface: #f2f2f2; --gm3-sys-color-inverse-on-surface-rgb: 242,242,242; --gm3-sys-color-inverse-primary: #a8c7fa; --gm3-sys-color-inverse-primary-rgb: 168,199,250; --gm3-sys-color-inverse-surface: #303030; --gm3-sys-color-inverse-surface-rgb: 48,48,48; --gm3-sys-color-on-background: #1f1f1f; --gm3-sys-color-on-background-rgb: 31,31,31; --gm3-sys-color-on-error: #fff; --gm3-sys-color-on-error-rgb: 255,255,255; --gm3-sys-color-on-error-container: #410e0b; --gm3-sys-color-on-error-container-rgb: 65,14,11; --gm3-sys-color-on-primary: #fff; --gm3-sys-color-on-primary-rgb: 255,255,255; --gm3-sys-color-on-primary-container: #041e49; --gm3-sys-color-on-primary-container-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed: #041e49; --gm3-sys-color-on-primary-fixed-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed-variant: #0842a0; --gm3-sys-color-on-primary-fixed-variant-rgb: 8,66,160; --gm3-sys-color-on-secondary: #fff; --gm3-sys-color-on-secondary-rgb: 255,255,255; --gm3-sys-color-on-secondary-container: #001d35; --gm3-sys-color-on-secondary-container-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed: #001d35; --gm3-sys-color-on-secondary-fixed-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed-variant: #004a77; --gm3-sys-color-on-secondary-fixed-variant-rgb: 0,74,119; --gm3-sys-color-on-surface: #1f1f1f; --gm3-sys-color-on-surface-rgb: 31,31,31; --gm3-sys-color-on-surface-variant: #444746; --gm3-sys-color-on-surface-variant-rgb: 68,71,70; --gm3-sys-color-on-tertiary: #fff; --gm3-sys-color-on-tertiary-rgb: 255,255,255; --gm3-sys-color-on-tertiary-container: #072711; --gm3-sys-color-on-tertiary-container-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed: #072711; --gm3-sys-color-on-tertiary-fixed-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed-variant: #0f5223; --gm3-sys-color-on-tertiary-fixed-variant-rgb: 15,82,35; --gm3-sys-color-outline: #747775; --gm3-sys-color-outline-rgb: 116,119,117; --gm3-sys-color-outline-variant: #c4c7c5; --gm3-sys-color-outline-variant-rgb: 196,199,197; --gm3-sys-color-primary: #0b57d0; --gm3-sys-color-primary-rgb: 11,87,208; --gm3-sys-color-primary-container: #d3e3fd; --gm3-sys-color-primary-container-rgb: 211,227,253; --gm3-sys-color-primary-fixed: #d3e3fd; --gm3-sys-color-primary-fixed-rgb: 211,227,253; --gm3-sys-color-primary-fixed-dim: #a8c7fa; --gm3-sys-color-primary-fixed-dim-rgb: 168,199,250; --gm3-sys-color-scrim: #000; --gm3-sys-color-scrim-rgb: 0,0,0; --gm3-sys-color-secondary: #00639b; --gm3-sys-color-secondary-rgb: 0,99,155; --gm3-sys-color-secondary-container: #c2e7ff; --gm3-sys-color-secondary-container-rgb: 194,231,255; --gm3-sys-color-secondary-fixed: #c2e7ff; --gm3-sys-color-secondary-fixed-rgb: 194,231,255; --gm3-sys-color-secondary-fixed-dim: #7fcfff; --gm3-sys-color-secondary-fixed-dim-rgb: 127,207,255; --gm3-sys-color-shadow: #000; --gm3-sys-color-shadow-rgb: 0,0,0; --gm3-sys-color-surface: #fff; --gm3-sys-color-surface-rgb: 255,255,255; --gm3-sys-color-surface-bright: #fff; --gm3-sys-color-surface-bright-rgb: 255,255,255; --gm3-sys-color-surface-container: #f0f4f9; --gm3-sys-color-surface-container-rgb: 240,244,249; --gm3-sys-color-surface-container-high: #e9eef6; --gm3-sys-color-surface-container-high-rgb: 233,238,246; --gm3-sys-color-surface-container-highest: #dde3ea; --gm3-sys-color-surface-container-highest-rgb: 221,227,234; --gm3-sys-color-surface-container-low: #f8fafd; --gm3-sys-color-surface-container-low-rgb: 248,250,253; --gm3-sys-color-surface-container-lowest: #fff; --gm3-sys-color-surface-container-lowest-rgb: 255,255,255; --gm3-sys-color-surface-dim: #d3dbe5; --gm3-sys-color-surface-dim-rgb: 211,219,229; --gm3-sys-color-surface-tint: #6991d6; --gm3-sys-color-surface-tint-rgb: 105,145,214; --gm3-sys-color-surface-variant: #e1e3e1; --gm3-sys-color-surface-variant-rgb: 225,227,225; --gm3-sys-color-tertiary: #146c2e; --gm3-sys-color-tertiary-rgb: 20,108,46; --gm3-sys-color-tertiary-container: #c4eed0; --gm3-sys-color-tertiary-container-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed: #c4eed0; --gm3-sys-color-tertiary-fixed-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed-dim: #6dd58c; --gm3-sys-color-tertiary-fixed-dim-rgb: 109,213,140; }

.XV0XSd.LgGVmb { --dt-background: rgb(32,33,36); --dt-on-background: rgb(232,234,237); --dt-on-background-secondary: rgb(154,160,166); --dt-outline: rgb(95,99,104); --dt-outline-variant: rgb(189,193,198); --dt-on-disabled: rgba(232,234,237,0.38); --dt-disabled: rgba(232,234,237,0.12); --dt-inverse-on-surface: rgb(60,64,67); --dt-inverse-surface: rgb(241,243,244); --dt-on-surface-secondary: rgb(154,160,166); --dt-on-surface-variant: rgb(154,160,166); --dt-on-surface: rgb(232,234,237); --dt-surface-tint: rgb(60,64,67); --dt-surface-variant: rgb(60,64,67); --dt-surface1: rgb(32,33,36); --dt-surface1-shadow: 0 1px 2px 0 rgba(0,0,0,0.3),0 1px 3px 1px rgba(0,0,0,0.15); --dt-surface2: rgb(32,33,36); --dt-surface2-shadow: 0 1px 2px 0 rgba(0,0,0,0.3),0 2px 6px 2px rgba(0,0,0,0.15); --dt-surface3: #36373a; --dt-surface3-shadow: 0 1px 3px 0 rgba(0,0,0,0.3),0 4px 8px 3px rgba(0,0,0,0.15); --dt-surface4: rgb(32,33,36); --dt-surface4-shadow: 0 2px 3px 0 rgba(0,0,0,0.3),0 6px 10px 4px rgba(0,0,0,0.15); --dt-surface5: rgb(32,33,36); --dt-surface5-shadow: 0 4px 4px 0 rgba(0,0,0,0.3),0 8px 12px 6px rgba(0,0,0,0.15); --dt-surface: rgb(32,33,36); --dt-scrim: rgba(32,33,36,0.87); --dt-scrim-2x: rgb(241,243,244); --dt-on-primary-container: rgb(210,227,252); --dt-on-primary: rgb(32,33,36); --dt-primary-action-state-layer: rgb(138,180,248); --dt-primary-action-stateful: rgb(174,203,250); --dt-primary-action: rgb(138,180,248); --dt-primary-container-icon: rgb(210,227,252); --dt-primary-container-link: rgb(210,227,252); --dt-primary-container: #394457; --dt-primary-icon: rgb(32,33,36); --dt-primary-link: rgb(32,33,36); --dt-primary-outline: rgb(138,180,248); --dt-primary: rgb(138,180,248); --dt-on-secondary-container: rgb(241,243,244); --dt-on-secondary: rgb(218,220,224); --dt-secondary-action-state-layer: rgb(218,220,224); --dt-secondary-action-stateful: rgb(232,234,237); --dt-secondary-action: rgb(218,220,224); --dt-secondary-container-icon: rgb(241,243,244); --dt-secondary-container-link: rgb(241,243,244); --dt-secondary-container: #4d4e51; --dt-secondary-icon: rgb(218,220,224); --dt-secondary-link: rgb(218,220,224); --dt-secondary-outline: rgb(218,220,224); --dt-secondary: rgb(32,33,36); --dt-on-tertiary-container: rgb(206,234,214); --dt-on-tertiary: rgb(32,33,36); --dt-tertiary-action-state-layer: rgb(129,201,149); --dt-tertiary-action-stateful: rgb(168,218,181); --dt-tertiary-action: rgb(129,201,149); --dt-tertiary-container-icon: rgb(206,234,214); --dt-tertiary-container-link: rgb(206,234,214); --dt-tertiary-container: #37493f; --dt-tertiary-icon: rgb(32,33,36); --dt-tertiary-link: rgb(32,33,36); --dt-tertiary-outline: rgb(129,201,149); --dt-tertiary: rgb(129,201,149); --dt-on-neutral-container: rgb(232,234,237); --dt-on-neutral: rgb(32,33,36); --dt-neutral-action-state-layer: rgb(232,234,237); --dt-neutral-action-stateful: #fff; --dt-neutral-action: rgb(232,234,237); --dt-neutral-container-icon: rgb(232,234,237); --dt-neutral-container-link: rgb(174,203,250); --dt-neutral-container: rgb(60,64,67); --dt-neutral-icon: rgb(32,33,36); --dt-neutral-link: rgb(32,33,36); --dt-neutral-outline: rgb(232,234,237); --dt-neutral: rgb(232,234,237); --dt-error-action-state-layer: rgb(242,139,130); --dt-error-action-stateful: rgb(246,174,169); --dt-error-action: rgb(242,139,130); --dt-error-container-icon: rgb(250,210,207); --dt-error-container-link: rgb(250,210,207); --dt-error-container: #523a3b; --dt-error-icon: rgb(32,33,36); --dt-error-link: rgb(32,33,36); --dt-error-outline: rgb(242,139,130); --dt-error: rgb(242,139,130); --dt-on-error-container: rgb(250,210,207); --dt-on-error: rgb(32,33,36); --dt-on-warning-container: rgb(254,239,195); --dt-on-warning: rgb(32,33,36); --dt-warning-action-state-layer: rgb(253,214,99); --dt-warning-action-stateful: rgb(253,226,147); --dt-warning-action: rgb(253,214,99); --dt-warning-container-icon: rgb(254,239,195); --dt-warning-container-link: rgb(254,239,195); --dt-warning-container: #554c33; --dt-warning-icon: rgb(32,33,36); --dt-warning-link: rgb(32,33,36); --dt-warning-outline: rgb(253,214,99); --dt-warning: rgb(253,214,99); --gm3-sys-color-background: #1f1f1f; --gm3-sys-color-background-rgb: 31,31,31; --gm3-sys-color-error: #f2b8b5; --gm3-sys-color-error-rgb: 242,184,181; --gm3-sys-color-error-container: #8c1d18; --gm3-sys-color-error-container-rgb: 140,29,24; --gm3-sys-color-inverse-on-surface: #303030; --gm3-sys-color-inverse-on-surface-rgb: 48,48,48; --gm3-sys-color-inverse-primary: #0b57d0; --gm3-sys-color-inverse-primary-rgb: 11,87,208; --gm3-sys-color-inverse-surface: #e3e3e3; --gm3-sys-color-inverse-surface-rgb: 227,227,227; --gm3-sys-color-on-background: #e3e3e3; --gm3-sys-color-on-background-rgb: 227,227,227; --gm3-sys-color-on-error: #601410; --gm3-sys-color-on-error-rgb: 96,20,16; --gm3-sys-color-on-error-container: #f9dedc; --gm3-sys-color-on-error-container-rgb: 249,222,220; --gm3-sys-color-on-primary: #062e6f; --gm3-sys-color-on-primary-rgb: 6,46,111; --gm3-sys-color-on-primary-container: #d3e3fd; --gm3-sys-color-on-primary-container-rgb: 211,227,253; --gm3-sys-color-on-primary-fixed: #041e49; --gm3-sys-color-on-primary-fixed-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed-variant: #0842a0; --gm3-sys-color-on-primary-fixed-variant-rgb: 8,66,160; --gm3-sys-color-on-secondary: #035; --gm3-sys-color-on-secondary-rgb: 0,51,85; --gm3-sys-color-on-secondary-container: #c2e7ff; --gm3-sys-color-on-secondary-container-rgb: 194,231,255; --gm3-sys-color-on-secondary-fixed: #001d35; --gm3-sys-color-on-secondary-fixed-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed-variant: #004a77; --gm3-sys-color-on-secondary-fixed-variant-rgb: 0,74,119; --gm3-sys-color-on-surface: #e3e3e3; --gm3-sys-color-on-surface-rgb: 227,227,227; --gm3-sys-color-on-surface-variant: #c4c7c5; --gm3-sys-color-on-surface-variant-rgb: 196,199,197; --gm3-sys-color-on-tertiary: #0a3818; --gm3-sys-color-on-tertiary-rgb: 10,56,24; --gm3-sys-color-on-tertiary-container: #c4eed0; --gm3-sys-color-on-tertiary-container-rgb: 196,238,208; --gm3-sys-color-on-tertiary-fixed: #072711; --gm3-sys-color-on-tertiary-fixed-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed-variant: #0f5223; --gm3-sys-color-on-tertiary-fixed-variant-rgb: 15,82,35; --gm3-sys-color-outline: #8e918f; --gm3-sys-color-outline-rgb: 142,145,143; --gm3-sys-color-outline-variant: #444746; --gm3-sys-color-outline-variant-rgb: 68,71,70; --gm3-sys-color-primary: #a8c7fa; --gm3-sys-color-primary-rgb: 168,199,250; --gm3-sys-color-primary-container: #0842a0; --gm3-sys-color-primary-container-rgb: 8,66,160; --gm3-sys-color-primary-fixed: #d3e3fd; --gm3-sys-color-primary-fixed-rgb: 211,227,253; --gm3-sys-color-primary-fixed-dim: #a8c7fa; --gm3-sys-color-primary-fixed-dim-rgb: 168,199,250; --gm3-sys-color-scrim: #000; --gm3-sys-color-scrim-rgb: 0,0,0; --gm3-sys-color-secondary: #7fcfff; --gm3-sys-color-secondary-rgb: 127,207,255; --gm3-sys-color-secondary-container: #004a77; --gm3-sys-color-secondary-container-rgb: 0,74,119; --gm3-sys-color-secondary-fixed: #c2e7ff; --gm3-sys-color-secondary-fixed-rgb: 194,231,255; --gm3-sys-color-secondary-fixed-dim: #7fcfff; --gm3-sys-color-secondary-fixed-dim-rgb: 127,207,255; --gm3-sys-color-shadow: #000; --gm3-sys-color-shadow-rgb: 0,0,0; --gm3-sys-color-surface: #1f1f1f; --gm3-sys-color-surface-rgb: 31,31,31; --gm3-sys-color-surface-bright: #37393b; --gm3-sys-color-surface-bright-rgb: 55,57,59; --gm3-sys-color-surface-container: #1e1f20; --gm3-sys-color-surface-container-rgb: 30,31,32; --gm3-sys-color-surface-container-high: #282a2c; --gm3-sys-color-surface-container-high-rgb: 40,42,44; --gm3-sys-color-surface-container-highest: #333537; --gm3-sys-color-surface-container-highest-rgb: 51,53,55; --gm3-sys-color-surface-container-low: #1b1b1b; --gm3-sys-color-surface-container-low-rgb: 27,27,27; --gm3-sys-color-surface-container-lowest: #0e0e0e; --gm3-sys-color-surface-container-lowest-rgb: 14,14,14; --gm3-sys-color-surface-dim: #131313; --gm3-sys-color-surface-dim-rgb: 19,19,19; --gm3-sys-color-surface-tint: #d1e1ff; --gm3-sys-color-surface-tint-rgb: 209,225,255; --gm3-sys-color-surface-variant: #444746; --gm3-sys-color-surface-variant-rgb: 68,71,70; --gm3-sys-color-tertiary: #6dd58c; --gm3-sys-color-tertiary-rgb: 109,213,140; --gm3-sys-color-tertiary-container: #0f5223; --gm3-sys-color-tertiary-container-rgb: 15,82,35; --gm3-sys-color-tertiary-fixed: #c4eed0; --gm3-sys-color-tertiary-fixed-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed-dim: #6dd58c; --gm3-sys-color-tertiary-fixed-dim-rgb: 109,213,140; }

.vhoiae.KkxPLb { --dt-on-background: #1F1F1F; --dt-on-background-secondary: #5E5E5E; --dt-background: #FFF; --dt-on-surface: #1F1F1F; --dt-inverse-surface: #303030; --dt-on-surface-secondary: #5E5E5E; --dt-on-surface-variant: #444746; --dt-surface-variant: #E3E3E3; --dt-inverse-on-surface: #F2F2F2; --dt-surface: #FFF; --dt-surface-tint: #6991d6; --dt-surface1: #f7f9fc; --dt-surface1-shadow: 0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12); --dt-surface2: #f2f6fc; --dt-surface2-shadow: 0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12); --dt-surface3: #edf2fc; --dt-surface3-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface4: #e8effb; --dt-surface4-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface5: #e2ecfb; --dt-surface5-shadow: 0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12); --dt-scrim: rgba(0,0,0,0.32); --dt-scrim-2x: rgba(0,0,0,0.64); --dt-on-primary-container: #041E49; --dt-primary-container-icon: #041E49; --dt-primary-container-link: #041E49; --dt-primary: #0B57D0; --dt-primary-action: #0B57D0; --dt-primary-action-stateful: #0B57D0; --dt-primary-outline: #0B57D0; --dt-primary-action-state-layer: #0B57D0; --dt-primary-container: #D3E3FD; --dt-on-primary: #FFF; --dt-primary-icon: #FFF; --dt-primary-link: #FFF; --dt-on-secondary-container: #001D35; --dt-secondary-container-icon: #001D35; --dt-secondary-container-link: #001D35; --dt-secondary: #00639B; --dt-secondary-action: #00639B; --dt-secondary-action-stateful: #00639B; --dt-secondary-outline: #00639B; --dt-secondary-action-state-layer: #00639B; --dt-secondary-container: #C2E7FF; --dt-on-secondary: #FFF; --dt-secondary-icon: #FFF; --dt-secondary-link: #FFF; --dt-on-tertiary-container: #072711; --dt-tertiary-container-icon: #072711; --dt-tertiary-container-link: #072711; --dt-tertiary: #146C2E; --dt-tertiary-action: #146C2E; --dt-tertiary-action-stateful: #146C2E; --dt-tertiary-outline: #146C2E; --dt-tertiary-action-state-layer: #146C2E; --dt-tertiary-container: #C4EED0; --dt-on-tertiary: #FFF; --dt-tertiary-icon: #FFF; --dt-tertiary-link: #FFF; --dt-on-neutral-container: #1F1F1F; --dt-neutral-container-icon: #1F1F1F; --dt-neutral-container-link: #1F1F1F; --dt-neutral: #474747; --dt-neutral-action: #1F1F1F; --dt-neutral-action-stateful: #1F1F1F; --dt-neutral-outline: #1F1F1F; --dt-neutral-action-state-layer: #1F1F1F; --dt-neutral-container: #E3E3E3; --dt-on-neutral: #FFF; --dt-neutral-icon: #FFF; --dt-neutral-link: #FFF; --dt-on-warning-container: #421F00; --dt-warning-container-icon: #421F00; --dt-warning-container-link: #421F00; --dt-warning: #F09D00; --dt-warning-action: #421F00; --dt-warning-action-stateful: #421F00; --dt-warning-outline: #421F00; --dt-warning-action-state-layer: #421F00; --dt-warning-container: #FFDF99; --dt-on-warning: #1F1F1F; --dt-warning-icon: #1F1F1F; --dt-warning-link: #1F1F1F; --dt-on-error-container: #410E0B; --dt-error-container-icon: #410E0B; --dt-error-container-link: #410E0B; --dt-error: #B3261E; --dt-error-action: #B3261E; --dt-error-action-stateful: #B3261E; --dt-error-outline: #B3261E; --dt-error-action-state-layer: #B3261E; --dt-error-container: #F9DEDC; --dt-on-error: #FFF; --dt-error-icon: #FFF; --dt-error-link: #FFF; --dt-disabled: rgba(31,31,31,0.12); --dt-on-disabled: rgba(31,31,31,0.38); --dt-outline: #747775; --dt-outline-variant: #C7C7C7; --gm3-sys-color-background: #fff; --gm3-sys-color-background-rgb: 255,255,255; --gm3-sys-color-error: #b3261e; --gm3-sys-color-error-rgb: 179,38,30; --gm3-sys-color-error-container: #f9dedc; --gm3-sys-color-error-container-rgb: 249,222,220; --gm3-sys-color-inverse-on-surface: #f2f2f2; --gm3-sys-color-inverse-on-surface-rgb: 242,242,242; --gm3-sys-color-inverse-primary: #a8c7fa; --gm3-sys-color-inverse-primary-rgb: 168,199,250; --gm3-sys-color-inverse-surface: #303030; --gm3-sys-color-inverse-surface-rgb: 48,48,48; --gm3-sys-color-on-background: #1f1f1f; --gm3-sys-color-on-background-rgb: 31,31,31; --gm3-sys-color-on-error: #fff; --gm3-sys-color-on-error-rgb: 255,255,255; --gm3-sys-color-on-error-container: #410e0b; --gm3-sys-color-on-error-container-rgb: 65,14,11; --gm3-sys-color-on-primary: #fff; --gm3-sys-color-on-primary-rgb: 255,255,255; --gm3-sys-color-on-primary-container: #041e49; --gm3-sys-color-on-primary-container-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed: #041e49; --gm3-sys-color-on-primary-fixed-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed-variant: #0842a0; --gm3-sys-color-on-primary-fixed-variant-rgb: 8,66,160; --gm3-sys-color-on-secondary: #fff; --gm3-sys-color-on-secondary-rgb: 255,255,255; --gm3-sys-color-on-secondary-container: #001d35; --gm3-sys-color-on-secondary-container-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed: #001d35; --gm3-sys-color-on-secondary-fixed-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed-variant: #004a77; --gm3-sys-color-on-secondary-fixed-variant-rgb: 0,74,119; --gm3-sys-color-on-surface: #1f1f1f; --gm3-sys-color-on-surface-rgb: 31,31,31; --gm3-sys-color-on-surface-variant: #444746; --gm3-sys-color-on-surface-variant-rgb: 68,71,70; --gm3-sys-color-on-tertiary: #fff; --gm3-sys-color-on-tertiary-rgb: 255,255,255; --gm3-sys-color-on-tertiary-container: #072711; --gm3-sys-color-on-tertiary-container-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed: #072711; --gm3-sys-color-on-tertiary-fixed-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed-variant: #0f5223; --gm3-sys-color-on-tertiary-fixed-variant-rgb: 15,82,35; --gm3-sys-color-outline: #747775; --gm3-sys-color-outline-rgb: 116,119,117; --gm3-sys-color-outline-variant: #c4c7c5; --gm3-sys-color-outline-variant-rgb: 196,199,197; --gm3-sys-color-primary: #0b57d0; --gm3-sys-color-primary-rgb: 11,87,208; --gm3-sys-color-primary-container: #d3e3fd; --gm3-sys-color-primary-container-rgb: 211,227,253; --gm3-sys-color-primary-fixed: #d3e3fd; --gm3-sys-color-primary-fixed-rgb: 211,227,253; --gm3-sys-color-primary-fixed-dim: #a8c7fa; --gm3-sys-color-primary-fixed-dim-rgb: 168,199,250; --gm3-sys-color-scrim: #000; --gm3-sys-color-scrim-rgb: 0,0,0; --gm3-sys-color-secondary: #00639b; --gm3-sys-color-secondary-rgb: 0,99,155; --gm3-sys-color-secondary-container: #c2e7ff; --gm3-sys-color-secondary-container-rgb: 194,231,255; --gm3-sys-color-secondary-fixed: #c2e7ff; --gm3-sys-color-secondary-fixed-rgb: 194,231,255; --gm3-sys-color-secondary-fixed-dim: #7fcfff; --gm3-sys-color-secondary-fixed-dim-rgb: 127,207,255; --gm3-sys-color-shadow: #000; --gm3-sys-color-shadow-rgb: 0,0,0; --gm3-sys-color-surface: #fff; --gm3-sys-color-surface-rgb: 255,255,255; --gm3-sys-color-surface-bright: #fff; --gm3-sys-color-surface-bright-rgb: 255,255,255; --gm3-sys-color-surface-container: #f0f4f9; --gm3-sys-color-surface-container-rgb: 240,244,249; --gm3-sys-color-surface-container-high: #e9eef6; --gm3-sys-color-surface-container-high-rgb: 233,238,246; --gm3-sys-color-surface-container-highest: #dde3ea; --gm3-sys-color-surface-container-highest-rgb: 221,227,234; --gm3-sys-color-surface-container-low: #f8fafd; --gm3-sys-color-surface-container-low-rgb: 248,250,253; --gm3-sys-color-surface-container-lowest: #fff; --gm3-sys-color-surface-container-lowest-rgb: 255,255,255; --gm3-sys-color-surface-dim: #d3dbe5; --gm3-sys-color-surface-dim-rgb: 211,219,229; --gm3-sys-color-surface-tint: #6991d6; --gm3-sys-color-surface-tint-rgb: 105,145,214; --gm3-sys-color-surface-variant: #e1e3e1; --gm3-sys-color-surface-variant-rgb: 225,227,225; --gm3-sys-color-tertiary: #146c2e; --gm3-sys-color-tertiary-rgb: 20,108,46; --gm3-sys-color-tertiary-container: #c4eed0; --gm3-sys-color-tertiary-container-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed: #c4eed0; --gm3-sys-color-tertiary-fixed-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed-dim: #6dd58c; --gm3-sys-color-tertiary-fixed-dim-rgb: 109,213,140; }

.vhoiae.LgGVmb { --dt-on-background: #E3E3E3; --dt-on-background-secondary: #ABABAB; --dt-background: #1F1F1F; --dt-on-surface: #E3E3E3; --dt-inverse-surface: #E3E3E3; --dt-on-surface-secondary: #ABABAB; --dt-on-surface-variant: #C4C7C5; --dt-surface-variant: #444746; --dt-inverse-on-surface: #303030; --dt-surface: #1F1F1F; --dt-surface-tint: #d1e1ff; --dt-surface1: #292a2d; --dt-surface1-shadow: 0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12); --dt-surface2: #2d2f33; --dt-surface2-shadow: 0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12); --dt-surface3: #31343a; --dt-surface3-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface4: #32363c; --dt-surface4-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface5: #353940; --dt-surface5-shadow: 0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12); --dt-scrim: rgba(0,0,0,0.32); --dt-scrim-2x: rgba(0,0,0,0.64); --dt-on-primary-container: #D3E3FD; --dt-primary-container-icon: #D3E3FD; --dt-primary-container-link: #D3E3FD; --dt-primary: #A8C7FA; --dt-primary-action: #A8C7FA; --dt-primary-action-stateful: #A8C7FA; --dt-primary-outline: #A8C7FA; --dt-primary-action-state-layer: #1B6EF3; --dt-primary-container: #0842A0; --dt-on-primary: #062E6F; --dt-primary-icon: #062E6F; --dt-primary-link: #062E6F; --dt-on-secondary-container: #C2E7FF; --dt-secondary-container-icon: #C2E7FF; --dt-secondary-container-link: #C2E7FF; --dt-secondary: #7FCFFF; --dt-secondary-action: #7FCFFF; --dt-secondary-action-stateful: #7FCFFF; --dt-secondary-outline: #7FCFFF; --dt-secondary-action-state-layer: #047DB7; --dt-secondary-container: #004A77; --dt-on-secondary: #035; --dt-secondary-icon: #035; --dt-secondary-link: #035; --dt-on-tertiary-container: #C4EED0; --dt-tertiary-container-icon: #C4EED0; --dt-tertiary-container-link: #C4EED0; --dt-tertiary: #6DD58C; --dt-tertiary-action: #6DD58C; --dt-tertiary-action-stateful: #6DD58C; --dt-tertiary-outline: #6DD58C; --dt-tertiary-action-state-layer: #198639; --dt-tertiary-container: #0F5223; --dt-on-tertiary: #0A3818; --dt-tertiary-icon: #0A3818; --dt-tertiary-link: #0A3818; --dt-on-neutral-container: #E3E3E3; --dt-neutral-container-icon: #E3E3E3; --dt-neutral-container-link: #E3E3E3; --dt-neutral: #ABABAB; --dt-neutral-action: #ABABAB; --dt-neutral-action-stateful: #ABABAB; --dt-neutral-outline: #ABABAB; --dt-neutral-action-state-layer: #ABABAB; --dt-neutral-container: #474747; --dt-on-neutral: #1F1F1F; --dt-neutral-icon: #ABABAB; --dt-neutral-link: #ABABAB; --dt-on-warning-container: #FFF0D1; --dt-warning-container-icon: #FFF0D1; --dt-warning-container-link: #FFF0D1; --dt-warning: #FFBB29; --dt-warning-action: #FFBB29; --dt-warning-action-stateful: #FFBB29; --dt-warning-outline: #FFF0D1; --dt-warning-action-state-layer: #FFBB29; --dt-warning-container: #562D00; --dt-on-warning: #1F1F1F; --dt-warning-icon: #421F00; --dt-warning-link: #421F00; --dt-on-error-container: #F9DEDC; --dt-error-container-icon: #F9DEDC; --dt-error-container-link: #F9DEDC; --dt-error: #F2B8B5; --dt-error-action: #F2B8B5; --dt-error-action-stateful: #F2B8B5; --dt-error-outline: #F2B8B5; --dt-error-action-state-layer: #DC362E; --dt-error-container: #8C1D18; --dt-on-error: #601410; --dt-error-icon: #601410; --dt-error-link: #601410; --dt-disabled: rgba(227,227,227,0.12); --dt-on-disabled: rgba(227,227,227,0.38); --dt-outline: #8E918F; --dt-outline-variant: #444746; --gm3-sys-color-background: #1f1f1f; --gm3-sys-color-background-rgb: 31,31,31; --gm3-sys-color-error: #f2b8b5; --gm3-sys-color-error-rgb: 242,184,181; --gm3-sys-color-error-container: #8c1d18; --gm3-sys-color-error-container-rgb: 140,29,24; --gm3-sys-color-inverse-on-surface: #303030; --gm3-sys-color-inverse-on-surface-rgb: 48,48,48; --gm3-sys-color-inverse-primary: #0b57d0; --gm3-sys-color-inverse-primary-rgb: 11,87,208; --gm3-sys-color-inverse-surface: #e3e3e3; --gm3-sys-color-inverse-surface-rgb: 227,227,227; --gm3-sys-color-on-background: #e3e3e3; --gm3-sys-color-on-background-rgb: 227,227,227; --gm3-sys-color-on-error: #601410; --gm3-sys-color-on-error-rgb: 96,20,16; --gm3-sys-color-on-error-container: #f9dedc; --gm3-sys-color-on-error-container-rgb: 249,222,220; --gm3-sys-color-on-primary: #062e6f; --gm3-sys-color-on-primary-rgb: 6,46,111; --gm3-sys-color-on-primary-container: #d3e3fd; --gm3-sys-color-on-primary-container-rgb: 211,227,253; --gm3-sys-color-on-primary-fixed: #041e49; --gm3-sys-color-on-primary-fixed-rgb: 4,30,73; --gm3-sys-color-on-primary-fixed-variant: #0842a0; --gm3-sys-color-on-primary-fixed-variant-rgb: 8,66,160; --gm3-sys-color-on-secondary: #035; --gm3-sys-color-on-secondary-rgb: 0,51,85; --gm3-sys-color-on-secondary-container: #c2e7ff; --gm3-sys-color-on-secondary-container-rgb: 194,231,255; --gm3-sys-color-on-secondary-fixed: #001d35; --gm3-sys-color-on-secondary-fixed-rgb: 0,29,53; --gm3-sys-color-on-secondary-fixed-variant: #004a77; --gm3-sys-color-on-secondary-fixed-variant-rgb: 0,74,119; --gm3-sys-color-on-surface: #e3e3e3; --gm3-sys-color-on-surface-rgb: 227,227,227; --gm3-sys-color-on-surface-variant: #c4c7c5; --gm3-sys-color-on-surface-variant-rgb: 196,199,197; --gm3-sys-color-on-tertiary: #0a3818; --gm3-sys-color-on-tertiary-rgb: 10,56,24; --gm3-sys-color-on-tertiary-container: #c4eed0; --gm3-sys-color-on-tertiary-container-rgb: 196,238,208; --gm3-sys-color-on-tertiary-fixed: #072711; --gm3-sys-color-on-tertiary-fixed-rgb: 7,39,17; --gm3-sys-color-on-tertiary-fixed-variant: #0f5223; --gm3-sys-color-on-tertiary-fixed-variant-rgb: 15,82,35; --gm3-sys-color-outline: #8e918f; --gm3-sys-color-outline-rgb: 142,145,143; --gm3-sys-color-outline-variant: #444746; --gm3-sys-color-outline-variant-rgb: 68,71,70; --gm3-sys-color-primary: #a8c7fa; --gm3-sys-color-primary-rgb: 168,199,250; --gm3-sys-color-primary-container: #0842a0; --gm3-sys-color-primary-container-rgb: 8,66,160; --gm3-sys-color-primary-fixed: #d3e3fd; --gm3-sys-color-primary-fixed-rgb: 211,227,253; --gm3-sys-color-primary-fixed-dim: #a8c7fa; --gm3-sys-color-primary-fixed-dim-rgb: 168,199,250; --gm3-sys-color-scrim: #000; --gm3-sys-color-scrim-rgb: 0,0,0; --gm3-sys-color-secondary: #7fcfff; --gm3-sys-color-secondary-rgb: 127,207,255; --gm3-sys-color-secondary-container: #004a77; --gm3-sys-color-secondary-container-rgb: 0,74,119; --gm3-sys-color-secondary-fixed: #c2e7ff; --gm3-sys-color-secondary-fixed-rgb: 194,231,255; --gm3-sys-color-secondary-fixed-dim: #7fcfff; --gm3-sys-color-secondary-fixed-dim-rgb: 127,207,255; --gm3-sys-color-shadow: #000; --gm3-sys-color-shadow-rgb: 0,0,0; --gm3-sys-color-surface: #1f1f1f; --gm3-sys-color-surface-rgb: 31,31,31; --gm3-sys-color-surface-bright: #37393b; --gm3-sys-color-surface-bright-rgb: 55,57,59; --gm3-sys-color-surface-container: #1e1f20; --gm3-sys-color-surface-container-rgb: 30,31,32; --gm3-sys-color-surface-container-high: #282a2c; --gm3-sys-color-surface-container-high-rgb: 40,42,44; --gm3-sys-color-surface-container-highest: #333537; --gm3-sys-color-surface-container-highest-rgb: 51,53,55; --gm3-sys-color-surface-container-low: #1b1b1b; --gm3-sys-color-surface-container-low-rgb: 27,27,27; --gm3-sys-color-surface-container-lowest: #0e0e0e; --gm3-sys-color-surface-container-lowest-rgb: 14,14,14; --gm3-sys-color-surface-dim: #131313; --gm3-sys-color-surface-dim-rgb: 19,19,19; --gm3-sys-color-surface-tint: #d1e1ff; --gm3-sys-color-surface-tint-rgb: 209,225,255; --gm3-sys-color-surface-variant: #444746; --gm3-sys-color-surface-variant-rgb: 68,71,70; --gm3-sys-color-tertiary: #6dd58c; --gm3-sys-color-tertiary-rgb: 109,213,140; --gm3-sys-color-tertiary-container: #0f5223; --gm3-sys-color-tertiary-container-rgb: 15,82,35; --gm3-sys-color-tertiary-fixed: #c4eed0; --gm3-sys-color-tertiary-fixed-rgb: 196,238,208; --gm3-sys-color-tertiary-fixed-dim: #6dd58c; --gm3-sys-color-tertiary-fixed-dim-rgb: 109,213,140; }

.XV0XSd .yYWAMb.bvmRsc, .XV0XSd .dif24c.bvmRsc { --dt-background: rgb(32,33,36); --dt-on-background: rgb(232,234,237); --dt-on-background-secondary: rgb(154,160,166); --dt-outline: rgb(95,99,104); --dt-outline-variant: rgb(189,193,198); --dt-on-disabled: rgba(232,234,237,0.38); --dt-disabled: rgba(232,234,237,0.12); --dt-inverse-on-surface: rgb(60,64,67); --dt-inverse-surface: rgb(241,243,244); --dt-on-surface-secondary: rgb(154,160,166); --dt-on-surface-variant: rgb(154,160,166); --dt-on-surface: rgb(232,234,237); --dt-surface-tint: rgb(60,64,67); --dt-surface-variant: rgb(60,64,67); --dt-surface1: rgb(32,33,36); --dt-surface1-shadow: 0 1px 2px 0 rgba(0,0,0,0.3),0 1px 3px 1px rgba(0,0,0,0.15); --dt-surface2: rgb(32,33,36); --dt-surface2-shadow: 0 1px 2px 0 rgba(0,0,0,0.3),0 2px 6px 2px rgba(0,0,0,0.15); --dt-surface3: #36373a; --dt-surface3-shadow: 0 1px 3px 0 rgba(0,0,0,0.3),0 4px 8px 3px rgba(0,0,0,0.15); --dt-surface4: rgb(32,33,36); --dt-surface4-shadow: 0 2px 3px 0 rgba(0,0,0,0.3),0 6px 10px 4px rgba(0,0,0,0.15); --dt-surface5: rgb(32,33,36); --dt-surface5-shadow: 0 4px 4px 0 rgba(0,0,0,0.3),0 8px 12px 6px rgba(0,0,0,0.15); --dt-surface: rgb(32,33,36); --dt-scrim: rgba(32,33,36,0.87); --dt-scrim-2x: rgb(241,243,244); --dt-on-primary-container: rgb(210,227,252); --dt-on-primary: rgb(32,33,36); --dt-primary-action-state-layer: rgb(138,180,248); --dt-primary-action-stateful: rgb(174,203,250); --dt-primary-action: rgb(138,180,248); --dt-primary-container-icon: rgb(210,227,252); --dt-primary-container-link: rgb(210,227,252); --dt-primary-container: #394457; --dt-primary-icon: rgb(32,33,36); --dt-primary-link: rgb(32,33,36); --dt-primary-outline: rgb(138,180,248); --dt-primary: rgb(138,180,248); --dt-on-secondary-container: rgb(241,243,244); --dt-on-secondary: rgb(218,220,224); --dt-secondary-action-state-layer: rgb(218,220,224); --dt-secondary-action-stateful: rgb(232,234,237); --dt-secondary-action: rgb(218,220,224); --dt-secondary-container-icon: rgb(241,243,244); --dt-secondary-container-link: rgb(241,243,244); --dt-secondary-container: #4d4e51; --dt-secondary-icon: rgb(218,220,224); --dt-secondary-link: rgb(218,220,224); --dt-secondary-outline: rgb(218,220,224); --dt-secondary: rgb(32,33,36); --dt-on-tertiary-container: rgb(206,234,214); --dt-on-tertiary: rgb(32,33,36); --dt-tertiary-action-state-layer: rgb(129,201,149); --dt-tertiary-action-stateful: rgb(168,218,181); --dt-tertiary-action: rgb(129,201,149); --dt-tertiary-container-icon: rgb(206,234,214); --dt-tertiary-container-link: rgb(206,234,214); --dt-tertiary-container: #37493f; --dt-tertiary-icon: rgb(32,33,36); --dt-tertiary-link: rgb(32,33,36); --dt-tertiary-outline: rgb(129,201,149); --dt-tertiary: rgb(129,201,149); --dt-on-neutral-container: rgb(232,234,237); --dt-on-neutral: rgb(32,33,36); --dt-neutral-action-state-layer: rgb(232,234,237); --dt-neutral-action-stateful: #fff; --dt-neutral-action: rgb(232,234,237); --dt-neutral-container-icon: rgb(232,234,237); --dt-neutral-container-link: rgb(174,203,250); --dt-neutral-container: rgb(60,64,67); --dt-neutral-icon: rgb(32,33,36); --dt-neutral-link: rgb(32,33,36); --dt-neutral-outline: rgb(232,234,237); --dt-neutral: rgb(232,234,237); --dt-error-action-state-layer: rgb(242,139,130); --dt-error-action-stateful: rgb(246,174,169); --dt-error-action: rgb(242,139,130); --dt-error-container-icon: rgb(250,210,207); --dt-error-container-link: rgb(250,210,207); --dt-error-container: #523a3b; --dt-error-icon: rgb(32,33,36); --dt-error-link: rgb(32,33,36); --dt-error-outline: rgb(242,139,130); --dt-error: rgb(242,139,130); --dt-on-error-container: rgb(250,210,207); --dt-on-error: rgb(32,33,36); --dt-on-warning-container: rgb(254,239,195); --dt-on-warning: rgb(32,33,36); --dt-warning-action-state-layer: rgb(253,214,99); --dt-warning-action-stateful: rgb(253,226,147); --dt-warning-action: rgb(253,214,99); --dt-warning-container-icon: rgb(254,239,195); --dt-warning-container-link: rgb(254,239,195); --dt-warning-container: #554c33; --dt-warning-icon: rgb(32,33,36); --dt-warning-link: rgb(32,33,36); --dt-warning-outline: rgb(253,214,99); --dt-warning: rgb(253,214,99); }

.vhoiae .yYWAMb.bvmRsc, .vhoiae .dif24c.bvmRsc, .X9XeLb .yYWAMb.bvmRsc, .X9XeLb .dif24c.bvmRsc, .cWKK1c .yYWAMb.bvmRsc, .cWKK1c .dif24c.bvmRsc, .aJfoSc .yYWAMb.bvmRsc, .aJfoSc .dif24c.bvmRsc, .TOb6Ze .yYWAMb.bvmRsc, .TOb6Ze .dif24c.bvmRsc { --dt-on-background: #E3E3E3; --dt-on-background-secondary: #ABABAB; --dt-background: #1F1F1F; --dt-on-surface: #E3E3E3; --dt-inverse-surface: #E3E3E3; --dt-on-surface-secondary: #ABABAB; --dt-on-surface-variant: #C4C7C5; --dt-surface-variant: #444746; --dt-inverse-on-surface: #303030; --dt-surface: #1F1F1F; --dt-surface-tint: #d1e1ff; --dt-surface1: #292a2d; --dt-surface1-shadow: 0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12); --dt-surface2: #2d2f33; --dt-surface2-shadow: 0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12); --dt-surface3: #31343a; --dt-surface3-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface4: #32363c; --dt-surface4-shadow: 0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12); --dt-surface5: #353940; --dt-surface5-shadow: 0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12); --dt-scrim: rgba(0,0,0,0.32); --dt-scrim-2x: rgba(0,0,0,0.64); --dt-on-primary-container: #D3E3FD; --dt-primary-container-icon: #D3E3FD; --dt-primary-container-link: #D3E3FD; --dt-primary: #A8C7FA; --dt-primary-action: #A8C7FA; --dt-primary-action-stateful: #A8C7FA; --dt-primary-outline: #A8C7FA; --dt-primary-action-state-layer: #1B6EF3; --dt-primary-container: #0842A0; --dt-on-primary: #062E6F; --dt-primary-icon: #062E6F; --dt-primary-link: #062E6F; --dt-on-secondary-container: #C2E7FF; --dt-secondary-container-icon: #C2E7FF; --dt-secondary-container-link: #C2E7FF; --dt-secondary: #7FCFFF; --dt-secondary-action: #7FCFFF; --dt-secondary-action-stateful: #7FCFFF; --dt-secondary-outline: #7FCFFF; --dt-secondary-action-state-layer: #047DB7; --dt-secondary-container: #004A77; --dt-on-secondary: #035; --dt-secondary-icon: #035; --dt-secondary-link: #035; --dt-on-tertiary-container: #C4EED0; --dt-tertiary-container-icon: #C4EED0; --dt-tertiary-container-link: #C4EED0; --dt-tertiary: #6DD58C; --dt-tertiary-action: #6DD58C; --dt-tertiary-action-stateful: #6DD58C; --dt-tertiary-outline: #6DD58C; --dt-tertiary-action-state-layer: #198639; --dt-tertiary-container: #0F5223; --dt-on-tertiary: #0A3818; --dt-tertiary-icon: #0A3818; --dt-tertiary-link: #0A3818; --dt-on-neutral-container: #E3E3E3; --dt-neutral-container-icon: #E3E3E3; --dt-neutral-container-link: #E3E3E3; --dt-neutral: #ABABAB; --dt-neutral-action: #ABABAB; --dt-neutral-action-stateful: #ABABAB; --dt-neutral-outline: #ABABAB; --dt-neutral-action-state-layer: #ABABAB; --dt-neutral-container: #474747; --dt-on-neutral: #1F1F1F; --dt-neutral-icon: #ABABAB; --dt-neutral-link: #ABABAB; --dt-on-warning-container: #FFF0D1; --dt-warning-container-icon: #FFF0D1; --dt-warning-container-link: #FFF0D1; --dt-warning: #FFBB29; --dt-warning-action: #FFBB29; --dt-warning-action-stateful: #FFBB29; --dt-warning-outline: #FFF0D1; --dt-warning-action-state-layer: #FFBB29; --dt-warning-container: #562D00; --dt-on-warning: #1F1F1F; --dt-warning-icon: #421F00; --dt-warning-link: #421F00; --dt-on-error-container: #F9DEDC; --dt-error-container-icon: #F9DEDC; --dt-error-container-link: #F9DEDC; --dt-error: #F2B8B5; --dt-error-action: #F2B8B5; --dt-error-action-stateful: #F2B8B5; --dt-error-outline: #F2B8B5; --dt-error-action-state-layer: #DC362E; --dt-error-container: #8C1D18; --dt-on-error: #601410; --dt-error-icon: #601410; --dt-error-link: #601410; --dt-disabled: rgba(227,227,227,0.12); --dt-on-disabled: rgba(227,227,227,0.38); --dt-outline: #8E918F; --dt-outline-variant: #444746; }

.I1PgQd { box-sizing: border-box; padding: 0.5rem 1rem; width: 20rem; }

.ousvBd { -webkit-box-align: center; align-items: center; display: flex; margin-right: -0.5rem; }

.Zcp8g.vKmmhc { color: var(--dt-on-surface,#3c4043); font-size: 1.25rem; line-height: 1.25rem; margin-right: 0.3rem; }

.nCnYNd { font: var(--dt-title-small-font,500 .875rem/1.25rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-small-spacing,0.0178571429em); color: var(--dt-on-surface,#3c4043); -webkit-box-flex: 1; flex: 1 1 0%; }

.EafEFe { font: var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-large-spacing,0); margin-bottom: 0.75rem; }

.RQM9Gf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); color: var(--dt-on-surface,#3c4043); }

.EIsVy { display: flex; -webkit-box-pack: end; justify-content: flex-end; margin: 0px -0.25rem; }

.BjbK3c { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; background: var(--dt-surface2,#fff); border-radius: 0.5rem; position: relative; }

.BjbK3c::before { border: 1px solid transparent; border-radius: inherit; inset: 0px; content: ""; position: absolute; }

.kaZy8e, .cDqddf, .FfqPSe, .kAgEFc { fill: var(--dt-background,#fff); position: absolute; }

.kaZy8e, .FfqPSe { height: 1.0625rem; left: 50%; margin-left: -0.9375rem; width: 1.875rem; }

.kaZy8e { top: -1.0625rem; }

.FfqPSe { bottom: -1.0625rem; }

.cDqddf, .kAgEFc { height: 1.875rem; margin-top: -0.9375rem; top: 50%; width: 1.0625rem; }

.cDqddf { right: -1.0625rem; }

.kAgEFc { left: -1.0625rem; }

.ob9sLd { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-stretch: ; font-size: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-small-spacing,.025em); border-radius: 0.25rem; box-sizing: border-box; display: inline-block; font-weight: 500; height: 1.25rem; line-height: 1.25rem; overflow: hidden; padding: 0px 0.5rem; position: relative; text-overflow: ellipsis; white-space: nowrap; }

.ob9sLd::before { border: 1px solid transparent; border-radius: inherit; inset: 0px; content: ""; position: absolute; }

@media (forced-colors: active) {
  .ob9sLd::before { border-color: canvastext; }
}

@media (forced-colors: active) {
  .RCmsv { background-color: buttonface !important; }
  .RCmsv, .RCmsv::before { border-color: buttontext !important; }
  .RCmsv:disabled, .RCmsv.RDPZE, .RCmsv:disabled::before, .RCmsv.RDPZE::before { border-color: graytext !important; opacity: 1 !important; }
  .RCmsv.u3bW4e, .RCmsv:focus, .RCmsv:hover, .hp3b6d.u3bW4e, .hp3b6d:focus, .hp3b6d:hover { background-color: highlight !important; }
  .RCmsv.u3bW4e, .RCmsv:focus, .RCmsv:hover, .hp3b6d.u3bW4e, .hp3b6d:focus, .hp3b6d:hover, .RCmsv.u3bW4e::before, .RCmsv:focus::before, .RCmsv:hover::before, .hp3b6d.u3bW4e::before, .hp3b6d:focus::before, .hp3b6d:hover::before { border-color: highlighttext !important; outline-color: highlighttext !important; }
  .jbArdc, .jbArdc [viewbox] { forced-color-adjust: none; color: buttontext !important; fill: currentcolor !important; }
  .jbArdc:disabled, .jbArdc.RDPZE, .jbArdc:disabled [viewbox], .jbArdc.RDPZE [viewbox] { color: graytext !important; opacity: 1 !important; }
  .jbArdc.u3bW4e, .jbArdc:focus, .jbArdc:hover, .jbArdc.u3bW4e [viewbox], .jbArdc:focus [viewbox], .jbArdc:hover [viewbox] { color: highlighttext !important; }
  .Yz4sEb { background-color: field !important; border-color: fieldtext !important; }
  .Yz4sEb:disabled, .Yz4sEb.RDPZE { border-color: graytext !important; }
  .GyDQo { forced-color-adjust: none; color: fieldtext !important; fill: currentcolor !important; }
  .GyDQo:disabled, .GyDQo.RDPZE { color: graytext !important; opacity: 1 !important; }
  .GyDQo::-webkit-input-placeholder { color: graytext !important; opacity: 1 !important; }
  .GyDQo::placeholder { color: graytext !important; opacity: 1 !important; }
  .cNqOse { background-color: canvas !important; }
  .cNqOse.kUXOd { border-color: canvastext !important; border-style: solid !important; border-width: 1px !important; }
  .X0gZEc { forced-color-adjust: none; color: canvastext !important; fill: currentcolor !important; }
  .ObwPwb { background-color: highlight !important; }
  .rkFgee { forced-color-adjust: none; color: highlighttext !important; fill: currentcolor !important; }
  .uevTLb { forced-color-adjust: none; color: linktext !important; fill: currentcolor !important; }
  .uevTLb:active, .uevTLb.qs41qe { color: activetext !important; }
  .uevTLb:visited, .uevTLb.gxDgLe { color: visitedtext !important; }
}

.HB1eCd-HzV7m .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge .HB1eCd-Bz112c, .HB1eCd-HzV7m .EX2EHc-INgbqf-hxXJme-xl07Ob-LgbsSe .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .HB1eCd-Bz112c { height: 18px; width: 18px; margin: 1px 2px 2px 1px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531.svg"); }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531.svg"); }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); }

.HB1eCd-fuEl3d-n9v5ye .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c-haAclf { height: 13220px; position: absolute; width: 83px; }

.HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-RJLb9c-haAclf { opacity: 0.54; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-RJLb9c-haAclf, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-OMz1o, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-usbjsf, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-EgTfg, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-hDEnYe, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-I9GLp, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-nA1mMd, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-wlNA0d, .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-jSFuyb { opacity: 1; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge .HB1eCd-Bz112c { margin-top: 0px; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c::before { content: ""; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c { content: ""; }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-HzV7m.lUepf-nEeMgc .HB1eCd-Bz112c { margin: 4px; }

.HB1eCd-HzV7m .HB1eCd-QbdDtf-oKdM2c-Bz112c .RbRzK-Bz112c { margin: -1px 0px 0px -1px; }

.HB1eCd-Bz112c-sLO9V-rdwzAe { font-family: "Google Symbols"; height: 0px; position: absolute; overflow: hidden; width: 0px; z-index: -1; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-w7bdYb-iyXyEd { left: 0px; top: -9674px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Q4BLdf { left: 0px; top: -9014px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-jNm5if { left: -40px; top: -7146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-HB1eCd { left: 0px; top: -11530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-RFAvhb { left: 0px; top: -11838px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-a1e4Ad { left: 0px; top: -2826px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-iyXyEd { left: 0px; top: -11818px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-xJzy8c { left: 0px; top: -9164px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-wcotoc-ndfHFb { left: -40px; top: -1438px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-cGMI2b { left: -40px; top: -3060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-oXtfBe { left: -60px; top: -3060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-oXtfBe { left: -20px; top: -8792px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-LK5yu { left: -26px; top: -7890px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-qwU8Me { left: -20px; top: -12210px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-yIbDgf { left: 0px; top: -2356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-LK5yu { left: 0px; top: -6876px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-AipIyc { left: 0px; top: -4020px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-qwU8Me { left: 0px; top: -12506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-ma6Yeb { left: -42px; top: -8690px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-cGMI2b { left: -48px; top: -13172px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-oXtfBe { left: -26px; top: -7646px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-ma6Yeb { left: -40px; top: -3102px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XXCpLd-Bpn8Yb { left: -62px; top: -11344px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XXCpLd-Bpn8Yb-mlk5z { left: -40px; top: -2978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-OiiCO { left: -22px; top: -11304px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KmuGVc-MHYjYb { left: -52px; top: -10648px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MqcBrc-s4vhY { left: -42px; top: -8730px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-IyROMc-wlNA0d { left: -40px; top: -10466px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o { left: -26px; top: -10012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o-v3pZbf { left: -20px; top: -76px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o-MFS4be { left: 0px; top: -2958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XHgP6b-SDqDXe-iAqvw { left: -62px; top: -3472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XHgP6b-f4z2Dd-E4ZlWe { left: -60px; top: -5388px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-elBQIf { left: -62px; top: -4964px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-c8csvc { left: -20px; top: -3594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-K0TrJc { left: -62px; top: -12668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-HrRdod-yLHjwb { left: -62px; top: -9634px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-km6h5c { left: 0px; top: -4882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QLEXN { left: -42px; top: -1062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QLEXN-DKlKme { left: -42px; top: -5708px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-WPi0i-MR5Q1e { left: 0px; top: -4964px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MPu53c { left: -26px; top: -10222px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-OVkoRd-GEUYHe { left: -15px; top: -484px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JbbQac-Wxxdob { left: 0px; top: -7532px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TvD9Pc { left: 0px; top: -1084px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nyE0bc { left: -42px; top: -1230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-J5uZjd-edvN0e { left: -42px; top: -8770px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-DyVDA { left: 0px; top: -5166px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-DyVDA-mPlZac { left: 0px; top: -11346px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-N7Eqid-GMvhG { left: 0px; top: -608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-MCEKJb { left: -22px; top: -11654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bKkSne-obrOwb { left: -26px; top: -10182px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bN97Pc-jCCvxc { left: -42px; top: -3472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bMcfAe-pKrx3d-lbYRR { left: -26px; top: -1014px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QdThLb { left: -60px; top: -12820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-UkZFS { left: -62px; top: -11304px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xceQUb { left: -20px; top: -8536px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-VkLyEc-zM6fo { left: -20px; top: -5388px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-FuIHKe-R1gDOc-MR5Q1e { left: -40px; top: -6168px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Oo0NPd { left: 0px; top: -3100px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uG5Yqe-JPn0pf-DKlKme { left: -20px; top: -9932px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uG5Yqe-JPn0pf-BvBYQ { left: 0px; top: -5086px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nupQLb { left: -20px; top: -11530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nupQLb-Q4BLdf { left: 0px; top: -2482px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-cXXICe-x5cW0b { left: -42px; top: -8710px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn { left: 0px; top: -7512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn-MFS4be { left: -60px; top: -2114px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn-oq6NAc { left: 0px; top: -12210px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ndfHFb-aTv5jf { left: 0px; top: -4546px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-j4gsHd-hFsbo-bEDTcc-LkdAo { left: 0px; top: -4040px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DyVDA-D5MPn { left: -20px; top: -12360px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DyVDA-D5MPn-ImBhed { left: -26px; top: -8624px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xvr5H-i5vt6e { left: 0px; top: -3182px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wz3zdc { left: -62px; top: -1230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DJPBic-AFZkUd { left: -20px; top: -3684px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fHSeKd-LkdAo { left: -26px; top: -6230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-vgRlPd-XigvTc-rDoBzb { left: 0px; top: -1062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KoToPc { left: -40px; top: -8792px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KoToPc-DKlKme { left: -40px; top: -9932px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hdBvUb { left: 0px; top: -6654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PlOyMe-vOE8Lb-jCCvxc { left: 0px; top: -3532px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TZk80d-ZGNLv-I9GLp { left: -20px; top: -12918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TZk80d-jCCvxc { left: 0px; top: -6586px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-HTFGIc { left: 0px; top: -12002px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-bRSSXe { left: 0px; top: -2868px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-bRSSXe-Hyc8Sd { left: -20px; top: -2754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-jyrRxf-nUpftc { left: -20px; top: -1698px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-lCdvJf-bEDTcc-DARUcf { left: 0px; top: -10648px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-lCdvJf-BIr6Bc { left: -20px; top: -3882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-drxrmf-wcotoc-jirZld { left: -62px; top: -11798px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-AHmuwe-oXtfBe { left: -20px; top: -3102px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yEEHq { left: -20px; top: -6028px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yEEHq-x5cW0b { left: -62px; top: -8150px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-JNdkSc { left: 0px; top: -13074px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-JPn0pf { left: -34px; top: -5926px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-xSQTrd { left: 0px; top: -7444px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sLO9V-fmcmS-SxQuSe { left: -40px; top: -11738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xRdasc-oKdM2c-dJDgTb { left: 0px; top: -4422px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n9oEIb { left: -44px; top: -8812px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n9oEIb-SNIJTd { left: -42px; top: -1738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TBCoIc { left: 0px; top: -3122px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ObfsIf-KzxUkd { left: -42px; top: -12688px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ObfsIf-vhhrIe { left: -40px; top: -5514px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-tJHJj-yePe5c { left: -26px; top: -6520px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-h9d3hd { left: -60px; top: -1498px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ZYIfFd-fbudBf { left: -60px; top: -2774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ntN8G { left: 0px; top: -5648px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TIHSC-E8fGCc { left: -52px; top: -8878px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DKlKme-RWgCYc { left: 0px; top: -3320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DKlKme-YMi5E { left: -20px; top: -5608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xguqbd { left: 0px; top: -10668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-YRhSCb { left: 0px; top: -1564px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-YRhSCb-SIsrTd { left: -62px; top: -5660px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-nGOfy { left: -42px; top: -12042px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-nGOfy-SIsrTd { left: -22px; top: -10716px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Tswv1b { left: -20px; top: -10472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-kWbB0e-D5MPn { left: -20px; top: -3554px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-YPqjbf { left: 0px; top: -12400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rYk4U { left: -42px; top: -4712px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-c53jI-TBCoIc { left: -20px; top: -8858px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-O807Gb { left: -60px; top: -8858px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-LIMNJb { left: 0px; top: -320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-LIMNJb-AznF2e { left: 0px; top: -232px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc { left: -62px; top: -7512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-mSEUvf { left: -52px; top: -9118px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-QLEXN-VMPhoe { left: -62px; top: -6762px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-wwuYjd { left: -20px; top: -7126px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-yY4Wcc { left: -20px; top: -2114px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd { left: -60px; top: -3882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd-Q4BLdf { left: -62px; top: -3280px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd-Xhs9z { left: -62px; top: -5708px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Jn51gd { left: -40px; top: -8476px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Jn51gd-SIsrTd { left: 0px; top: -5388px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Rv62Se { left: -42px; top: -4628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pGuBYc-TvD9Pc { left: -62px; top: -6742px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pGuBYc-FNFY6c { left: -20px; top: -10758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-l4eHX-t02dhe { left: 0px; top: -8750px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JtB1fc { left: -52px; top: -7404px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xSh02c { left: -20px; top: -10506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-H1aTHf { left: -42px; top: -10310px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DUGJie-Q4BLdf { left: 0px; top: -3574px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-z5C9Gb-zcdHbf-BvBYQ { left: 0px; top: -4146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-x5cW0b-nKQ6qf-hgHJW { left: -40px; top: -4292px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-x5cW0b-nKQ6qf-yHKmmc { left: -42px; top: -7512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-h1U9Be { left: 0px; top: -7424px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RFnRab-MCEKJb { left: -60px; top: -9320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-b3rLgd-HzFBSb { left: -20px; top: -2336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Vgu1H-mKZypf { left: -22px; top: -1738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n5AaSd-u3Agqb { left: 0px; top: -1800px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PrY1nf-nQ1Faf { left: -60px; top: -9400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PrY1nf-nQ1Faf-MFS4be { left: -40px; top: -10958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pBztBd-dJfz0c-JZnCve { left: -40px; top: -12102px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-G84jIc { left: -62px; top: -3842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-FNFY6c-RmniWd-uJ3wk { left: -62px; top: -3662px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-LhcNjd { left: -22px; top: -12022px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-ij8cu { left: 0px; top: -5514px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-Lr2Z8d { left: 0px; top: -2436px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RF62N-nEeMgc-Ia7Qfc { left: 0px; top: -10472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KNM5Ef { left: -20px; top: -6210px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KNM5Ef-Q4BLdf { left: -40px; top: -212px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-g7W7Ed-qwU8Me-wcotoc-LK5yu { left: 0px; top: -170px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Ft5J4b { left: -62px; top: -4984px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Ft5J4b-di8rgd-Wxxdob { left: 0px; top: -9932px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-GEUYHe-JNdkSc { left: -26px; top: -7032px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Faem2b-cVFi4 { left: -48px; top: -8572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-iyXyEd { left: -48px; top: -1014px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-iyXyEd-g6cJHd { left: 0px; top: -11264px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nQ1Faf { left: -22px; top: -3202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nQ1Faf-Xhs9z { left: -26px; top: -9538px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xJzy8c-HiaYvf { left: -44px; top: -4400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xJzy8c-HiaYvf-O1htCb { left: 0px; top: -12420px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Jz7rA { left: 0px; top: -980px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-zSI2l-QLEXN { left: 0px; top: -6168px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n8nH7-jyrRxf { left: 0px; top: -9206px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jRmmHf-ibnC6b { left: -20px; top: -6676px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NziyQe-LkdAo { left: -52px; top: -6518px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TdyTDe { left: -20px; top: -5688px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TdyTDe-r9oPif { left: 0px; top: -9138px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-g3I98d { left: 0px; top: -2242px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-aIWppb-htvI8d { left: -46px; top: -5044px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EgTfg { left: -40px; top: -3554px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EgTfg-gS7Ybc { left: -40px; top: -2876px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PEFSMe { left: 0px; top: -9320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xXq91c-oQYOj { left: 0px; top: -4292px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Gpz5id { left: -40px; top: -8858px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uXLMpd { left: -60px; top: -8536px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qrlFte { left: -22px; top: -11674px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Iqlsrf { left: -58px; top: -6068px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-S9gUrf-HiaYvf { left: -60px; top: -10486px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-m3mY0d-Q4BLdf { left: 0px; top: -12380px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qwU8Me-rrhWne { left: 0px; top: -8792px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ReqAjb-qwU8Me-MnhZ9d { left: 0px; top: -8834px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ktSouf { left: -40px; top: -12820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NgtDm-YS35zb { left: -54px; top: -5004px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-O1htCb-NkyfNe { left: -20px; top: -11490px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EnFNjd-ryxqyc { left: -40px; top: -2814px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JPn0pf { left: 0px; top: -10248px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RFAvhb-AznF2e { left: -26px; top: -2502px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-if5aCc-sTBVle { left: -42px; top: -11674px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-luNtDf-s2ctBd { left: 0px; top: -13116px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-V5oUn { left: -20px; top: -2868px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb { left: -60px; top: -10506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb-e7aFhf { left: -20px; top: -1438px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb-uTrtOd { left: -40px; top: -2336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rvOPdc-RFnRab { left: 0px; top: -300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JK9eJ { left: 0px; top: -8496px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DIdRlc { left: -40px; top: -11510px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DIdRlc-nyE0bc { left: 0px; top: -8690px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hDEnYe-JaPV2b { left: -22px; top: -2548px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hDEnYe-nllRtd { left: 0px; top: -5668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-Q4BLdf-gvZm2b { left: -20px; top: -608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-ObfsIf-nUpftc { left: 0px; top: -8476px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-uaxL4e { left: -62px; top: -1130px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i2RYZ { left: 0px; top: -192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sTBVle-BvBYQ { left: -52px; top: -7424px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Yygnk { left: -42px; top: -11404px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Yygnk-Z5I80b { left: -26px; top: -7672px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-QLEXN { left: -60px; top: -6296px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-g6cJHd { left: -40px; top: -11550px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-AznF2e { left: -42px; top: -11654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-sAb8f { left: -60px; top: -3902px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-rrhWne-hgHJW { left: -20px; top: -5988px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-rrhWne-yHKmmc { left: -20px; top: -9952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-hgHJW { left: 0px; top: -5146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-tSZMSb { left: 0px; top: -3902px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-yHKmmc { left: -20px; top: -6190px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-BvBYQ-EbqdBd { left: -60px; top: -3080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EWK8Bb { left: -20px; top: -2958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RCfa3e { left: -62px; top: -252px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-L4Nn5e { left: -20px; top: -11940px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-e3BBL-yHKmmc-hFsbo { left: -20px; top: -11510px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Zj4Smb-Z5I80b-GMvhG { left: 0px; top: -1020px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NowJzb { left: 0px; top: -6316px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sfGayb { left: -42px; top: -11818px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MHYjYb-J6RZ7b { left: -40px; top: -8750px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-zf3vf { left: 0px; top: -3594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-dIxMhd-DyVDA-TIHSC { left: 0px; top: -6008px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-dIxMhd-iWMRLe-EnFNjd { left: 0px; top: -11570px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BvBYQ-nyE0bc { left: -46px; top: -12460px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nUpftc-kPTQic { left: -60px; top: -2436px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nUpftc-ti6hGc { left: -22px; top: -2896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qPaVXd-yHKmmc { left: 0px; top: -212px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PJVNOc-hYO5Oc { left: -42px; top: -8670px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-ltEGzf { left: 0px; top: -8858px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-RPzgNd { left: 0px; top: -4822px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-i8xkGf { left: -40px; top: -12230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nJjxad-bEDTcc { left: -58px; top: -5278px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-h30Snd-ovCUCd { left: -42px; top: -12002px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-h30Snd-ovCUCd-r9oPif { left: -46px; top: -9206px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb-ovCUCd { left: 0px; top: -340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ktSouf { left: -60px; top: -2978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PEFSMe { left: -60px; top: -12506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PEFSMe-E3DyYd { left: -20px; top: -1252px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb, .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-SIsrTd { left: -40px; top: -6028px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-E3DyYd, .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-SIsrTd-E3DyYd { left: -20px; top: -8670px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd, .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-SIsrTd { left: 0px; top: -6546px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-E3DyYd, .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-SIsrTd-E3DyYd { left: -58px; top: -2592px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc { left: 0px; top: -12820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc-r9oPif { left: -26px; top: -4080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-UkZFS { left: 0px; top: -11510px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b { left: -60px; top: -12860px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-OMz1o { left: 0px; top: -11408px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EgTfg, .HB1eCd-HzV7m .HB1eCd-Bz112c-usbjsf { left: -20px; top: -2436px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EgTfg-TLxrU { left: 0px; top: -11124px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hDEnYe { left: -60px; top: -9300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-I9GLp { left: 0px; top: -10268px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-I9GLp-JaPV2b { left: -60px; top: -6276px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd { left: -52px; top: -4754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jSFuyb { left: -40px; top: -9300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd-JaPV2b { left: 0px; top: -1458px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd-JaPV2b-r9oPif { left: -40px; top: -5682px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TFrYib { left: -40px; top: -11880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-oO2eQ { left: 0px; top: -2628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PJVNOc { left: 0px; top: -10758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-wlNA0d { left: 0px; top: -3040px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-wlNA0d { left: -20px; top: -7444px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jbwjpc-RvIlWb { left: -52px; top: -9834px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lcE6r-JLm1tf-YZ04zc-RvIlWb { left: -52px; top: -4566px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-N7Eqid-RvIlWb { left: 0px; top: -8218px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-Xhs9z-RvIlWb { left: 0px; top: -5900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vVQOP { left: -40px; top: -7356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-AV3gEe-Q4BLdf-XpSwdc { left: 0px; top: -10426px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf { left: -48px; top: -1034px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eFD6re { left: 0px; top: -6722px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-c8csvc { left: -20px; top: -668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-c8csvc-E3DyYd { left: 0px; top: -6632px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-O807Gb { left: -62px; top: -9786px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-O807Gb-E3DyYd { left: -22px; top: -11716px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-hxXJme { left: -40px; top: -1458px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-hxXJme-E3DyYd { left: 0px; top: -2528px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-LK5yu { left: -62px; top: -6830px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-LK5yu-E3DyYd { left: 0px; top: -9538px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-oXtfBe { left: -40px; top: -2958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-oXtfBe-E3DyYd { left: -20px; top: -2072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-qwU8Me { left: -20px; top: -2978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-qwU8Me-E3DyYd { left: -20px; top: -3512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-yIbDgf { left: -62px; top: -12918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-yIbDgf-E3DyYd { left: 0px; top: -11980px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-LK5yu { left: -48px; top: -1938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-oXtfBe { left: 0px; top: -7356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-qwU8Me { left: -52px; top: -11084px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-ma6Yeb { left: 0px; top: -7124px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-AipIyc { left: -20px; top: -8650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-cGMI2b { left: -60px; top: -9932px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uG5Yqe-JPn0pf-agdLee { left: 0px; top: -1872px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uG5Yqe-JPn0pf-o7abwc { left: -40px; top: -6190px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-ma6Yeb { left: 0px; top: -12572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-ma6Yeb-E3DyYd { left: 0px; top: -9054px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-AipIyc { left: 0px; top: -10938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-AipIyc-E3DyYd { left: 0px; top: -6402px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-cGMI2b { left: 0px; top: -1438px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-cGMI2b-E3DyYd { left: -26px; top: -7592px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H { left: -26px; top: -6588px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-E3DyYd { left: 0px; top: -4712px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-r9oPif { left: -48px; top: -1370px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Rv62Se-EXHrde-Ca4zAd { left: 0px; top: -6424px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv { left: 0px; top: -11758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-E3DyYd { left: -60px; top: -5470px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-r9oPif { left: -20px; top: -12400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Jn51gd-EXHrde-Ca4zAd { left: -22px; top: -2722px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld { left: -26px; top: -9482px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-E3DyYd { left: -20px; top: -6456px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc { left: 0px; top: -6742px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-E3DyYd { left: -46px; top: -6230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd { left: 0px; top: -1000px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-E3DyYd { left: -46px; top: -5064px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nyE0bc { left: -20px; top: -11798px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NowJzb { left: -62px; top: -1110px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NowJzb-E3DyYd { left: -36px; top: -170px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-yTCTk { left: -20px; top: -3534px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-I7wDP { left: -48px; top: -7772px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-I7wDP-r9oPif-T60B1 { left: 0px; top: -12460px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf { left: 0px; top: -10918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf-E3DyYd { left: -52px; top: -5900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf-r9oPif-gS7Ybc { left: -26px; top: -582px; }

.HB1eCd-HzV7m .EX2EHc-Bz112c-LSk3jc-BHsdwc { left: 0px; top: -10114px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QBLLGd { left: -55px; top: -5112px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-weuhHc-E3DyYd { left: -48px; top: -9254px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-FXrc0c { left: 0px; top: -6190px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-wZVHld-V67aGc { left: -52px; top: -6696px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tJiF1e { left: 0px; top: -3362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MYFTse { left: -22px; top: -6916px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-di8rgd-hxXJme { left: 0px; top: -6230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-edvN0e-hxXJme { left: -60px; top: -2918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-edvN0e-hxXJme-E3DyYd { left: -26px; top: -3018px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-hxXJme { left: -40px; top: -3902px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-rTEl { left: -20px; top: -11694px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-SX9D7d-E3DyYd { left: 0px; top: -3842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf { left: -40px; top: -6722px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-r9oPif { left: 0px; top: -7572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-nUpftc-ZdbLkb { left: -60px; top: -9054px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-eKpHRd-BPrWId-r9oPif { left: -46px; top: -11224px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if { left: -42px; top: -9676px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-jNm5if-E3DyYd { left: -52px; top: -8594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e { left: -20px; top: -3122px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-E3DyYd { left: -48px; top: -13094px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-AHUcCb { left: -60px; top: -4060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-E3Uge { left: -20px; top: -1498px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-Qs3R8d-E3DyYd { left: -60px; top: -7356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-uPjwvb-ZdbLkb { left: -42px; top: -12572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-jNm5if { left: -20px; top: -2242px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-jNm5if-r9oPif { left: 0px; top: -2774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-yHKmmc-r9oPif { left: -48px; top: -12184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-yHKmmc-yaNpec { left: 0px; top: -9744px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-hgHJW-yaNpec { left: 0px; top: -7336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QLEXN { left: -20px; top: -3162px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-QLEXN-E3DyYd { left: -42px; top: -6916px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QLEXN-r9oPif { left: -48px; top: -7572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-SIsrTd { left: -22px; top: -8770px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-SIsrTd-E3DyYd { left: -52px; top: -3382px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-SIsrTd { left: -62px; top: -11384px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-SIsrTd-E3DyYd { left: -60px; top: -11940px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-SIsrTd { left: -60px; top: -8750px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-SIsrTd-E3DyYd { left: -20px; top: -9744px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-SIsrTd { left: 0px; top: -4842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-SIsrTd-E3DyYd { left: -26px; top: -9254px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-SIsrTd { left: 0px; top: -5106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-SIsrTd-E3DyYd { left: -42px; top: -1252px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-i3jM8c { left: -22px; top: -9676px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-i3jM8c-E3DyYd { left: -60px; top: -9952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-SIsrTd { left: -40px; top: -11530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-SIsrTd-E3DyYd { left: -60px; top: -6168px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vOE8Lb-SIsrTd { left: 0px; top: -11244px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vOE8Lb-SIsrTd-E3DyYd { left: -44px; top: -10978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf { left: 0px; top: -862px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LQY1ye { left: -62px; top: -11858px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zjQX3e { left: -62px; top: -4692px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i2RYZ { left: -60px; top: -3554px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i2RYZ-E3DyYd { left: 0px; top: -11284px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JbbQac-TCl01b { left: -20px; top: -5514px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd { left: -40px; top: -1498px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-E3DyYd { left: 0px; top: -7166px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-dJfz0c-JZnCve { left: -42px; top: -3300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-dJfz0c-JZnCve-r9oPif { left: -56px; top: -5952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-HLvlvd { left: -42px; top: -11304px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-purZT { left: 0px; top: -668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-SdkFre { left: 0px; top: -1758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RF62N-Wxxdob { left: -20px; top: -11738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RF62N-Wxxdob-E3DyYd { left: -20px; top: -11570px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf { left: -52px; top: -7444px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL { left: -40px; top: -12062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL-SIsrTd { left: 0px; top: -2754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DARUcf-LhcNjd { left: -22px; top: -12042px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DARUcf-LhcNjd-r9oPif { left: -22px; top: -13120px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc { left: 0px; top: -1658px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd { left: -62px; top: -9766px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yHKmmc { left: 0px; top: -1892px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hgHJW { left: 0px; top: -5608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-DARUcf { left: -48px; top: -9718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xvr5H { left: -20px; top: -3492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vgRlPd { left: -48px; top: -1918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vgRlPd-r9oPif { left: 0px; top: -2046px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DKlKme-RWgCYc { left: 0px; top: -3684px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DKlKme-RWgCYc-r9oPif { left: 0px; top: -3778px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-oXtfBe-VBrcT { left: -22px; top: -4712px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-oXtfBe-cGMI2b-VBrcT { left: -60px; top: -2754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-LK5yu-VBrcT { left: -20px; top: -628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-qwU8Me-VBrcT { left: -42px; top: -2072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mQXP-r9oPif { left: -40px; top: -5634px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-CtVXDf-r08add-BKD3ld-cXXICe-VBrcT { left: -26px; top: -9472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-NkyfNe { left: -62px; top: -10248px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-NkyfNe-E3DyYd { left: -46px; top: -1084px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-qwU8Me { left: 0px; top: -7146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-qwU8Me-E3DyYd { left: -22px; top: -4942px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-LK5yu { left: 0px; top: -6856px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-LK5yu-E3DyYd { left: -48px; top: -1820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-ma6Yeb { left: -26px; top: -9906px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-ma6Yeb-E3DyYd { left: -22px; top: -11980px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-cGMI2b { left: 0px; top: -12918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-cGMI2b-E3DyYd { left: -52px; top: -4774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-sfSLhd { left: 0px; top: -4166px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-sfSLhd-E3DyYd { left: -48px; top: -9608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-EcYfVc { left: -20px; top: -9184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-EcYfVc-E3DyYd { left: -48px; top: -8432px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-tSZMSb { left: 0px; top: -11694px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-tSZMSb-E3DyYd { left: -20px; top: -10526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-DKlKme { left: -62px; top: -8770px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-DKlKme-E3DyYd { left: 0px; top: -6498px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-BvBYQ { left: -62px; top: -11878px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-BvBYQ-E3DyYd { left: 0px; top: -6916px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xSh02c { left: -20px; top: -2826px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf { left: -40px; top: -12210px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd { left: -26px; top: -12460px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pXHOFf { left: 0px; top: -5024px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pXHOFf-MFS4be { left: -20px; top: -4060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-s2ctBd { left: -26px; top: -556px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-s2ctBd-E3DyYd { left: -52px; top: -2154px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-NUaK6d { left: -20px; top: -1892px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-PoC6nf { left: -46px; top: -7890px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-PoC6nf-i5vt6e { left: -44px; top: -7910px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e { left: -20px; top: -12526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e-ZmdkE { left: -22px; top: -1718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e-QDgCrf { left: 0px; top: -5628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-Hyc8Sd { left: 0px; top: -9184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb { left: -52px; top: -9492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-LkdAo-r9oPif { left: 0px; top: -7844px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-hJDwNd { left: 0px; top: -38px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-hJDwNd-sM5MNb { width: 36px; height: 36px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-a4fUwd { left: -60px; top: -8792px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-a4fUwd-SIsrTd { left: -60px; top: -11510px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-z5C9Gb { left: -26px; top: -3804px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-z5C9Gb-SIsrTd { left: 0px; top: -11880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-UlV2sd-OMz1o { left: -42px; top: -1758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-uPjwvb { left: -26px; top: -9808px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-h0Nkge-uPjwvb-r9oPif { left: 0px; top: -3804px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qrlFte-uPjwvb-r9oPif { left: -48px; top: -9880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd { left: -48px; top: -12142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-E3Uge { left: 0px; top: -11798px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-NkyfNe { left: -48px; top: -1418px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PJVNOc-hYO5Oc { left: 0px; top: -12082px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-PvhD9 { left: 0px; top: -2938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ij8cu-r9oPif { left: -52px; top: -11592px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd { left: -20px; top: -11960px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe { left: 0px; top: -5688px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe-HLvlvd { left: -60px; top: -8476px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-O0r3Gd { left: -40px; top: -1564px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-O0r3Gd-u0pjoe-r9oPif-Qhstab { left: -20px; top: -4822px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zM6fo { left: -22px; top: -1758px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8 { left: -40px; top: -6362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8-E3Uge { left: 0px; top: -7870px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pmuK7 { left: 0px; top: -7104px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-fZiSAe { left: -42px; top: -9786px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pX1iqf-kPTQic { left: -40px; top: -6830px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-SNIJTd-kPTQic { left: 0px; top: -5126px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-DyVDA { left: 0px; top: -11940px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-DyVDA-ImBhed { left: -26px; top: -4800px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-nUpftc { left: -60px; top: -2336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd { left: -26px; top: -9144px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-VCkuzd-TLxrU { left: 0px; top: -6456px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-VCkuzd-HLvlvd { left: -42px; top: -12918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-iyXyEd-TLxrU { left: 0px; top: -10958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-iyXyEd-JH1xTd-TLxrU { left: -20px; top: -3142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd-htvI8d-HLvlvd { left: -26px; top: -6628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc { left: -22px; top: -12688px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lbYRR { left: 0px; top: -842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d { left: -42px; top: -10072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G84jIc { left: 0px; top: -7012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-V67aGc-S8vSze { left: 0px; top: -4692px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pKrx3d-SxQuSe { left: -60px; top: -10526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xXq91c { left: 0px; top: -7378px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-T3yXSc { left: 0px; top: -12840px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-BvBYQ-kolMJb { left: -42px; top: -12708px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LK5yu-kqOKYb { left: -62px; top: -8670px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qwU8Me-kqOKYb { left: 0px; top: -12062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LK5yu-kqOKYb-kolMJb { left: -20px; top: -9320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qwU8Me-kqOKYb-kolMJb { left: 0px; top: -12800px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf { left: -20px; top: -4292px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-x5cW0b { left: -20px; top: -3902px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DltcQc-CCJ0ld { left: -22px; top: -4732px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NMrWyd-s3Bhse { left: -52px; top: -8218px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hj4D6d-vJ7A6b { left: -60px; top: -1658px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-bEDTcc-E3DyYd { left: -20px; top: -1062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-m9bMae { left: -26px; top: -8078px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-yY4Wcc { left: -62px; top: -4628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nupQLb { left: 0px; top: -6676px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MrxDPd-jyrRxf { left: 0px; top: -1110px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hDEnYe-jkpPIb { left: 0px; top: -11920px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-Q9HdGd { left: -20px; top: -4106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QbShld { left: 0px; top: -6382px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zcdHbf { left: 0px; top: -12122px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sJY2Bf-bVEB4e { left: -40px; top: -3492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf { left: 0px; top: -6566px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-OiiCO { left: -40px; top: -3882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-r9oPif { left: 0px; top: -530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-u0pjoe-u2z5K { left: -42px; top: -2180px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sKFHqe { left: -20px; top: -13074px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sKFHqe-SIsrTd { left: -20px; top: -6168px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NBDE7b { left: -46px; top: -3822px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod { left: -60px; top: -2794px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-CBeBSd-EFlEBf { left: 0px; top: -9634px; }

.HB1eCd-HzV7m .HB1eCd-VgwJlc-xTMeO { left: -20px; top: -4964px; }

.HB1eCd-HzV7m .HB1eCd-VgwJlc-FNFY6c { left: -60px; top: -608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc { left: -20px; top: -4984px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc-r9oPif { left: -48px; top: -2998px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ud7fr { left: -20px; top: -11880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-R1s0ee-uDEFge-yaNpec { left: 0px; top: -816px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ud7fr-r9oPif { left: -20px; top: -10622px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-v3pZbf { left: -62px; top: -3300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-aVTXAb { left: -40px; top: -2754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sI3MNd { left: -52px; top: -12754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed { left: -52px; top: -10710px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-E3DyYd { left: -52px; top: -10688px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc-JaPV2b { left: -26px; top: -2998px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-aVTXAb-v3pZbf { left: -60px; top: -9360px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc { left: -62px; top: -10132px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c { left: -62px; top: -10288px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c-rTEl { left: -40px; top: -4106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-rTEl { left: -26px; top: -6608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-rTEl { left: 0px; top: -4902px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl { left: -40px; top: -4146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl-E3DyYd { left: -52px; top: -9564px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl-r9oPif { left: -48px; top: -7078px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GCYh9b-rTEl { left: -46px; top: -816px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-skjTt-rTEl { left: -40px; top: -9320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-rTEl { left: 0px; top: -3080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ihIZgd-rTEl { left: -26px; top: -7572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-r9oPif { left: -56px; top: -6382px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-fmcmS-eEGnhe { left: -22px; top: -6402px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-IT5dJd { left: 0px; top: -7798px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-IT5dJd-HLvlvd { left: -62px; top: -4822px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-Xhs9z { left: -26px; top: -4334px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-nGOfy { left: -52px; top: -12552px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-nGOfy-E3DyYd { left: 0px; top: -1348px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-YRhSCb { left: 0px; top: -10526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-YRhSCb-E3DyYd { left: 0px; top: -4922px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-HLvlvd { left: -52px; top: -11042px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-di8rgd-YwNhXd { left: -22px; top: -4692px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QdThLb { left: -42px; top: -10052px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QdThLb-E3DyYd { left: 0px; top: -2846px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nllRtd-g6cJHd { left: -42px; top: -4250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sLO9V-SxQuSe { left: -52px; top: -10668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf-HiaYvf { left: -20px; top: -10918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf-HiaYvf-E3DyYd { left: 0px; top: -9608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YIAiIb-rDoBzb { left: -60px; top: -4106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Fq92xe-mU4ghb { left: -22px; top: -9634px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yUKnc { left: 0px; top: -2978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-RPzgNd { left: -56px; top: -6408px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-i8xkGf { left: 0px; top: -2134px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-ltEGzf { left: 0px; top: -2092px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-b58pU { left: -62px; top: -11818px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nllRtd-a4fUwd { left: -20px; top: -11346px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-HLvlvd { left: -26px; top: -3228px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-HLvlvd-SIsrTd { left: 0px; top: -9808px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-h9d3hd { left: -20px; top: -5470px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sn54Q-nllRtd { left: -52px; top: -8918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eNZ9Nb { left: -26px; top: -7614px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-r9oPif { left: -46px; top: -9906px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-JaPV2b { left: -60px; top: -2876px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-JaPV2b-nNtqDd { left: -40px; top: -2794px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-nllRtd { left: -20px; top: -1544px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-HLvlvd { left: -22px; top: -11324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-OpAKde-QLEXN { left: -20px; top: -12062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-OpAKde-QLEXN-HLvlvd { left: -22px; top: -4922px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-bEDTcc { left: -22px; top: -7166px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc { left: -60px; top: -3100px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc-i5vt6e-J9pn5c-r9oPif { left: -52px; top: -4592px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW { left: -44px; top: -11980px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW-i5vt6e-J9pn5c-r9oPif { left: 0px; top: -9560px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jsmBPd-GMvhG { left: -26px; top: -2482px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KsV2dd { left: -62px; top: -10052px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb { left: 0px; top: -6048px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-B1neQd-TCl01b { left: -40px; top: -9184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-UmQjBf { left: -20px; top: -6742px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-QLEXN { left: -58px; top: -5298px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-to915 { left: -26px; top: -9558px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-qwU8Me-IFdKyd-HLvlvd-r9oPif { left: -52px; top: -10896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-to915-SIsrTd { left: -46px; top: -2396px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc { left: -52px; top: -10156px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-E3DyYd { left: -20px; top: -10312px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-r9oPif { left: -52px; top: -10176px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-N2TEqe { left: -42px; top: -9766px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ZMv3u-QLEXN { left: 0px; top: -12898px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ZMv3u-QLEXN-i5vt6e-r9oPif { left: -26px; top: -6336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-dJDgTb-QLEXN { left: -62px; top: -10072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-dJDgTb-QLEXN-i5vt6e-r9oPif { left: -26px; top: -6562px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QLEXN { left: -62px; top: -11324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QLEXN-r9oPif { left: -44px; top: -4922px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN { left: -22px; top: -1230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN-i5vt6e { height: 18px; left: 0px; top: -10288px; width: 18px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN-i5vt6e-r9oPif { left: -48px; top: -3340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Cs2axe-vhhrIe { left: -40px; top: -2222px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-J6RZ7b { left: -62px; top: -1062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S { left: -40px; top: -3574px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S-r9oPif { left: 0px; top: -1912px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S-i5vt6e { left: -40px; top: -1544px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-RWgCYc-yY4Wcc { left: -62px; top: -12938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-RWgCYc-yY4Wcc-BHsdwc { left: 0px; top: -6126px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-uiYelc { left: -40px; top: -10486px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NBDE7b-JaPV2b { left: -42px; top: -12668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-yHKmmc { left: 0px; top: -9472px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-yHKmmc-E3DyYd { left: -40px; top: -6872px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-hgHJW { left: 0px; top: -9300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-hgHJW-E3DyYd { left: -20px; top: -3996px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-lm6F6 { left: -22px; top: -2528px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-lm6F6-E3DyYd { left: 0px; top: -10716px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-X808Kb { left: -52px; top: -1872px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-X808Kb-E3DyYd { left: -22px; top: -4670px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-BvBYQ { left: 0px; top: -12526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-BvBYQ-E3DyYd { left: -42px; top: -5492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-tSZMSb { left: -40px; top: -2774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-tSZMSb-E3DyYd { left: 0px; top: -1718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q0hgme-mSEUvf { left: -40px; top: -5388px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-jyrRxf { left: 0px; top: -8454px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-nKQ6qf { left: 0px; top: -6896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RPzgNd-vfifzc-RxYbNe { left: 0px; top: -8650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-E8fGCc { left: 0px; top: -5988px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-t6UvL { left: -20px; top: -9300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-cGMI2b { left: -26px; top: -10202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-LK5yu { left: -52px; top: -6564px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-qwU8Me { left: 0px; top: -11224px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-ma6Yeb { left: -26px; top: -8412px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-tsZdxf-HLvlvd { left: -62px; top: -1718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-T3iPGc-r9oPif { left: -40px; top: -3142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-zf3vf { left: 0px; top: -12102px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-zf3vf-r9oPif { left: 0px; top: -2456px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Jz7rA { left: -56px; top: -6428px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Jz7rA-r9oPif { left: -26px; top: -7818px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LIMNJb { left: -26px; top: -4754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KsV2dd-HLvlvd { left: -40px; top: -13074px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-QIk5de-OWB6Me-EFlEBf { left: -40px; top: -76px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ntN8G { left: -40px; top: -2918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RCfa3e { left: -62px; top: -7552px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd-HLvlvd { left: -42px; top: -11384px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd { left: -42px; top: -11344px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-bBybbf { left: -60px; top: -5514px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf { left: 0px; top: -7490px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-Xhs9z { left: -20px; top: -9014px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qPaVXd-yHKmmc { left: -62px; top: -10112px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qPaVXd-yHKmmc-MFS4be-u2z5K { left: -22px; top: -12860px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-km6h5c { left: 0px; top: -7058px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-km6h5c-i5vt6e-r9oPif { left: -26px; top: -10156px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-n8nH7-jyrRxf { left: 0px; top: -3142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-n8nH7-jyrRxf { left: 0px; top: -6362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c-QUIbkc-HLvlvd-GoS4Be { left: 0px; top: -9340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-feLNVc { left: 0px; top: -4126px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-feLNVc-r9oPif { left: -40px; top: -274px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe { left: -20px; top: -12102px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic { left: -62px; top: -300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-drxrmf-DKlKme { left: -42px; top: -4020px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-drxrmf-BvBYQ { left: -22px; top: -1396px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ReqAjb-XaHFse { left: 0px; top: -12308px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb { left: -52px; top: -11104px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-E3Uge { left: -20px; top: -9034px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-ZdbLkb { left: -22px; top: -11000px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-uPjwvb-ZdbLkb { left: 0px; top: -3340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g3I98d { left: -20px; top: -12840px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-elBQIf { left: -62px; top: -11694px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vVewSc { left: -22px; top: -3842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-bMcfAe { left: -20px; top: -192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-oPu43-E3DyYd { left: -60px; top: -1478px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-oPu43-r9oPif { left: -26px; top: -9502px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-uDEFge-to915-r9oPif-oVleVe { left: -22px; top: -1370px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-i5vt6e-E3DyYd { left: -20px; top: -5492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-i5vt6e-r9oPif { left: 0px; top: -934px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e { left: -26px; top: -1934px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e-E3DyYd { left: -42px; top: -6654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e-r9oPif { left: 0px; top: -9420px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-i5vt6e-r9oPif { left: 0px; top: -8598px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-i5vt6e-E3DyYd { left: -20px; top: -8244px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-MFS4be-r9oPif-aOn1pf { left: 0px; top: -5044px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-i5vt6e-E3DyYd { left: -20px; top: -9206px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-i5vt6e-r9oPif { left: -22px; top: -13146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf-i5vt6e-E3DyYd { left: 0px; top: -2722px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf-i5vt6e-r9oPif { left: 0px; top: -7032px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ihIZgd-i5vt6e-E3DyYd { left: 0px; top: -8324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HTJzpc-i5vt6e-E3DyYd { left: 0px; top: -4250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-w7bdYb { left: -26px; top: -8192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GEUYHe-r9oPif { left: -26px; top: -12328px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL-HLvlvd { left: -42px; top: -10132px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe { left: -40px; top: -9972px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe { left: -20px; top: -212px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif { left: 0px; top: -7078px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif-v3pZbf { left: -34px; top: -9340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif-HLvlvd { left: 0px; top: -8412px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-uPjwvb-RvIlWb { left: -20px; top: -1084px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-CwllA-E3DyYd { left: 0px; top: -3280px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-E3Uge-E3DyYd { left: 0px; top: -13198px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-r9oPif { left: 0px; top: -4336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-HLvlvd-r9oPif { left: -26px; top: -5336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-r9oPif { left: -22px; top: -3340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-HLvlvd-r9oPif { left: -52px; top: -10202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-hgHJW-r9oPif { left: 0px; top: -582px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-yHKmmc-r9oPif { left: -46px; top: -1518px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-r9oPif { left: -48px; top: -7464px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-E3Uge-r9oPif { left: 0px; top: -9854px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nEeMgc { left: -22px; top: -11284px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RFAvhb-jyrRxf-r9oPif { left: 0px; top: -4374px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-r9oPif { left: -20px; top: -11224px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-auswjd-r9oPif { left: -52px; top: -6606px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-Xhs9z-r9oPif { left: 0px; top: -252px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-E3DyYd { left: 0px; top: -10978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ { left: -60px; top: -9380px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ-E3DyYd { left: 0px; top: -12668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ-RvIlWb { left: -52px; top: -9092px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-ibnC6b { left: -20px; top: -8750px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XHoCPb-r9oPif-CwllA { left: -44px; top: -8832px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-jbwjpc { left: 0px; top: -3512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-N7Eqid-W3lGp { left: -58px; top: -12250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-H8nU8b-W3lGp { left: -16px; top: -5004px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-RPzgNd-vfifzc-RxYbNe-W3lGp { left: -26px; top: -7910px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-r9oPif { left: -26px; top: -6696px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-kODWGd { left: 0px; top: -1172px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-yEEHq { left: 0px; top: -8670px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ge6pde-LkdAo-QG5zS { left: 0px; top: -8516px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pI3EI { left: -40px; top: -12360px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e { left: -20px; top: -3040px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-nQ1Faf-E3DyYd { left: 0px; top: -5804px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-E3DyYd { left: 0px; top: -2896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-HLvlvd { left: -40px; top: -9992px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-nUpftc-YuD1xf { left: -20px; top: -300px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-nUpftc-YuD1xf-IT5dJd-iBxYy-hxXJme-AHe6Kc { left: -22px; top: -6382px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf { left: -40px; top: -2938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf-IT5dJd-iBxYy-hxXJme-AHe6Kc { left: 0px; top: -12754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf-mPlZac { left: -22px; top: -12668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc { left: 0px; top: -11738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc-HLvlvd { left: 0px; top: -8150px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc-FNFY6c { left: -22px; top: -4400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { left: 0px; top: -10506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY-r9oPif { left: 0px; top: -7672px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-p2N3pf-r9oPif { left: -22px; top: -12184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-N7Eqid { left: -22px; top: -4628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-DcLNVc-r9oPif { left: 0px; top: -9092px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-hgHJW { left: -34px; top: -5004px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-yHKmmc { left: -62px; top: -10268px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c-E3Uge { left: -52px; top: -11022px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ij8cu-E3Uge { left: -62px; top: -3594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc-uFfGwd { left: -52px; top: -6498px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JNdkSc { left: -42px; top: -6126px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-iMG1U-E3Uge { left: 0px; top: -12486px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc-c4YZDc-r9oPif-HLvlvd { left: 0px; top: -6696px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ugYG9-c4YZDc { left: -20px; top: -11264px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ugYG9-c4YZDc-r9oPif-HLvlvd { left: 0px; top: -7646px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc-r9oPif-HLvlvd { left: -42px; top: -2528px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc-r9oPif-HLvlvd { left: 0px; top: -7890px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk { left: -60px; top: -3574px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-rYk4U { left: 0px; top: -3492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-oScmOd { left: -20px; top: -4848px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-oScmOd { left: 0px; top: -12142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-oScmOd { left: 0px; top: -5216px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-FMvwCe-oScmOd { left: -20px; top: -320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-FMvwCe-oScmOd { left: 0px; top: -12938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-FMvwCe-oScmOd { left: 0px; top: -2180px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-u2z5K { left: -22px; top: -9054px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-u2z5K { left: -20px; top: -11900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-u2z5K { left: 0px; top: -6276px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-QymXn-u2z5K { left: -26px; top: 0px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-JeMQb { left: 0px; top: -10548px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-JeMQb { left: 0px; top: -1274px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-JeMQb { left: 0px; top: -2648px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-JeMQb { left: 0px; top: -12980px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-JeMQb { left: 0px; top: -7188px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-fmcmS { left: -40px; top: -608px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-fmcmS { left: -42px; top: -10290px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-fmcmS { left: -42px; top: -9634px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-fmcmS { left: -20px; top: -5106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-SfQLQb-fmcmS { left: -60px; top: -7012px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-SfQLQb-fmcmS { left: -22px; top: -3452px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-fmcmS { left: -52px; top: -6632px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-fmcmS { left: -40px; top: -1658px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-fmcmS { left: -22px; top: -12002px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-fmcmS { left: 0px; top: -5258px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-LK5yu-Ysl7Fe { left: 0px; top: -8350px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-oXtfBe-Ysl7Fe { left: 0px; top: -4566px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-qwU8Me-Ysl7Fe { left: 0px; top: -11592px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-LK5yu-Ysl7Fe { left: -26px; top: -952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-Ysl7Fe { left: 0px; top: -8878px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-qwU8Me-Ysl7Fe { left: 0px; top: -5408px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-LK5yu-Ysl7Fe { left: -26px; top: -4500px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-oXtfBe-Ysl7Fe { left: 0px; top: -11048px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-qwU8Me-Ysl7Fe { left: -26px; top: -11428px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qknJed-AFZkUd { left: 0px; top: -4060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-qknJed-AFZkUd-hJDwNd { left: -62px; top: -3642px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JLm1tf-DJPBic-AFZkUd-W3lGp-TLxrU { left: -46px; top: -3804px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RFnRab-r9oPif { left: 0px; top: -10690px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd { left: -60px; top: -3040px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc { left: -42px; top: -3452px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-aOn1pf { left: -20px; top: -4272px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-VqDHhd { left: -62px; top: -10092px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc { left: -62px; top: -1150px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc-E3DyYd { left: -20px; top: -3080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me { left: -20px; top: -6722px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-aOn1pf { left: -20px; top: -7146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd-r9oPif { left: -48px; top: -1892px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-r9oPif { left: 0px; top: -2998px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-r9oPif-aOn1pf { left: 0px; top: -2502px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-r9oPif-VqDHhd { left: -52px; top: -4080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc-r9oPif { left: -22px; top: -13094px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-r9oPif { left: -46px; top: -11124px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-r9oPif-aOn1pf { left: 0px; top: -556px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb { left: 0px; top: -2072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-JaPV2b { left: 0px; top: -960px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-r9oPif { left: -55px; top: -5086px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-r9oPif-gS7Ybc { left: 0px; top: -6830px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG { left: 0px; top: -9280px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-r9oPif { left: -52px; top: -1846px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-MFS4be-ETmUib { left: 0px; top: -5470px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-SeBwEf { left: -26px; top: -7844px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-SeBwEf-r9oPif { left: -20px; top: -4166px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b { left: -20px; top: -1478px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-GjlSrc { left: 0px; top: -648px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-V7AMae { left: -20px; top: -12820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-CwllA { left: 0px; top: -1544px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ONu0F { left: 0px; top: -8556px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-r9oPif { left: 0px; top: -2800px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-i5vt6e-TY4T7c { left: -20px; top: -4650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-E3DyYd { left: -20px; top: -12572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-r9oPif { left: -26px; top: -12728px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-r9oPif { left: -22px; top: -3616px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d { left: -42px; top: -6456px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-r9oPif { left: 0px; top: -882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq { left: -62px; top: -7532px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-VtOx3e { left: 0px; top: -1678px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-MFS4be { left: 0px; top: -76px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-Q4BLdf { left: -20px; top: -8476px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-r9oPif { left: 0px; top: -10012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-di8rgd-r9oPif { left: -42px; top: -3202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-Hjleke-r9oPif { left: 0px; top: -5336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-iOyk4d-r9oPif { left: 0px; top: -4520px; }

.HB1eCd-HzV7m .HB1eCd-bVEB4e { left: -20px; top: -12230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nGOfy-Dy7EIf { left: -52px; top: -2046px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YRhSCb-Dy7EIf { left: -42px; top: -3996px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ryxqyc-vUjI9d-hxGuWb { left: 0px; top: -484px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ryxqyc-pDPzzb-hxGuWb { left: -40px; top: -5086px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-muPwQb { left: -35px; top: -484px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-x5cW0b { left: 0px; top: -11778px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-ma6Yeb-LK5yu { left: 0px; top: -5926px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-ma6Yeb-qwU8Me { left: 0px; top: -3452px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-vbnc8b { left: 0px; top: -4106px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-vbnc8b-r9oPif { left: -52px; top: -9538px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-r9oPif { left: -20px; top: -9228px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-r9oPif-HLvlvd { left: 0px; top: -9906px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-Qs3R8d-RvIlWb { left: -52px; top: -556px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-Qs3R8d-RvIlWb { left: -40px; top: -5608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-uPjwvb-RvIlWb { left: -52px; top: -9808px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-uPjwvb-RvIlWb { left: 0px; top: -12546px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-r9oPif { left: 0px; top: -10156px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-LSK72c-r9oPif { left: -26px; top: -7378px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-LrF0Pc-r9oPif { left: 0px; top: -4080px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-r9oPif { left: -26px; top: -8594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-tcqZEf-r9oPif { left: -46px; top: -7844px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-LrF0Pc-r9oPif { left: 0px; top: -2376px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YxWbQd-r9oPif { left: 0px; top: -908px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YxWbQd { left: -20px; top: -3320px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb { left: 0px; top: -4650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-ZdbLkb { left: 0px; top: -10896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-uPjwvb-ZdbLkb { left: 0px; top: -7464px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-QLEXN-ZdbLkb { left: -52px; top: -7820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-wvGCSb-LoDsGd-jJ3Q2c-Q7Syqe-r9oPif { left: 0px; top: -11428px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8-HLvlvd { left: -20px; top: -8130px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RxTQ8e-oq6NAc { left: -26px; top: -4374px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Y5dbrb-r9oPif { left: -26px; top: -12546px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KNM5Ef { left: -40px; top: -3684px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue { left: -26px; top: -5044px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue-r9oPif { left: 0px; top: -9254px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue-RAze1d-r9oPif { left: -22px; top: -7464px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-r9oPif-aOn1pf { left: 0px; top: -7398px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-clhnwb { left: -40px; top: -8536px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e4raY { left: 0px; top: -9952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-rYk4U { left: -40px; top: -7012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vOBb1e { left: -40px; top: -2436px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-smkJ3e { left: 0px; top: -12360px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YJL97b { left: -62px; top: -4250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YJL97b-r9oPif { left: -46px; top: -8192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-tSZMSb { left: -40px; top: -9952px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-m3mY0d-RbRzK { left: -44px; top: -9696px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-M1QMZb-fmcmS { left: -20px; top: -10958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c { left: -20px; top: -4146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb { left: -58px; top: -170px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-W3lGp { left: 0px; top: -6762px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-E3DyYd { left: -40px; top: -5874px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-r9oPif { left: -46px; top: -12400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-Wz3zdc-Z7HxEc-r9oPif-T60B1 { left: -26px; top: -8218px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-Wz3zdc-Z7HxEc-LrF0Pc-r9oPif { left: 0px; top: -5186px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-hWJfub-yHKmmc-r9oPif-T60B1 { left: -26px; top: -9118px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-oSWire { left: -40px; top: -5470px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe { left: -22px; top: -4250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-E3DyYd { left: -22px; top: -9696px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-r9oPif { left: -22px; top: -13172px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-Qs3R8d-RvIlWb { left: 0px; top: -10202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Faem2b-cVFi4-r9oPif-mPlZac { left: 0px; top: -5362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-V67aGc-i5vt6e { left: 0px; top: -6028px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c-C2S4ob { left: 0px; top: -2114px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd-G0jgYd-r9oPif { left: 0px; top: -6250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-n6j7Re { left: -40px; top: -232px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uaxL4e-n6j7Re { left: 0px; top: -1478px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-h976Ve { left: -46px; top: -7646px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-ctOWCc-r9oPif { left: -48px; top: -9420px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eizL8e-Vgu1H-r9oPif { left: -26px; top: -2154px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-npMLoc-r9oPif { left: -20px; top: -11124px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop { left: 0px; top: -4272px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-E3DyYd { left: 0px; top: -4314px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-r9oPif { left: -46px; top: -10622px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-SIsrTd { left: -20px; top: -6048px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-SIsrTd-E3DyYd { left: 0px; top: -8812px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe { left: 0px; top: -9654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-HLvlvd { left: -26px; top: -4314px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-zYyPae { left: 0px; top: -13136px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-GjlSrc { left: 0px; top: -2222px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-V7AMae { left: -20px; top: -7424px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-CwllA { left: -42px; top: -11324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-gNuiOc-r9oPif { left: -26px; top: -9092px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-gNuiOc-HLvlvd-r9oPif { left: -46px; top: -836px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed { left: -20px; top: -2094px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-r9oPif { left: 0px; top: -7598px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-clPPge-r9oPif { left: -26px; top: -5900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-clPPge-E3DyYd { left: -40px; top: -3594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-r9oPif { left: -48px; top: -13142px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-u5Azmc { left: -20px; top: -6362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-LBRlSe { left: 0px; top: -12440px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GnPzId { left: -20px; top: -232px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-xZDoyc-MJ0UK { left: -40px; top: -12506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-a2ItGd { left: 0px; top: -13054px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-wWDucd { left: -40px; top: -4650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GEUYHe { left: -20px; top: -7012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-WX1Rmf { left: -20px; top: -3060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-c6tfMc { left: 0px; top: -3554px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e3uGsb { left: -40px; top: -2114px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-e3uGsb-C2NXRc { left: -40px; top: -10446px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc { left: -26px; top: -9854px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-I3TTMc { left: -60px; top: -9340px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-I3TTMc-nQ1Faf { left: -20px; top: -1658px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-r9oPif { left: -52px; top: -10922px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-E3DyYd { left: -20px; top: -5708px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-nUpftc-mG3Az-r9oPif { left: -52px; top: -11618px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-bstyQc { left: -20px; top: -2938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-u5Azmc-r9oPif { left: 0px; top: -9512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-LBRlSe-r9oPif { left: -52px; top: -12774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GnPzId-r9oPif { left: 0px; top: -11022px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-xZDoyc-MJ0UK-r9oPif { left: 0px; top: -8192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-a2ItGd-r9oPif { left: -22px; top: -1820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-wWDucd-r9oPif { left: 0px; top: -3228px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GEUYHe-r9oPif { left: -52px; top: -10870px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-WX1Rmf-r9oPif { left: -46px; top: -8624px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-c6tfMc-r9oPif { left: -48px; top: -13116px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-hauLI-ETmUib { left: 0px; top: -11490px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-hauLI-r9oPif-ETmUib { left: -46px; top: -7672px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JEruSd-ETmUib { left: 0px; top: -5492px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd-r9oPif { left: -42px; top: -8324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-JEruSd-r9oPif-ETmUib { left: 0px; top: -9972px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-r9oPif { left: 0px; top: -8078px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-E3DyYd { left: 0px; top: -11654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-uPjwvb-E3DyYd { left: -42px; top: -1778px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-E3DyYd-t24pnf { left: 0px; top: -13094px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic-mlKF6d-kRWtF { left: 0px; top: -10052px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic-LkdAo { left: -22px; top: -8324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-YjoMNe { left: -34px; top: -5968px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YjoMNe-IFdKyd { left: -20px; top: -842px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-YjoMNe-HLvlvd { left: 0px; top: -3882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-V5oUn { left: -20px; top: -8692px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H { left: -26px; top: -2416px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-h976Ve-r9oPif { left: -48px; top: -530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-YjoMNe-IFdKyd-r9oPif { left: -35px; top: -504px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-h976Ve { left: 0px; top: -1252px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-muPwQb-LSK72c-r9oPif { left: 0px; top: -8572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd { left: -48px; top: -5362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-LkdAo { left: 0px; top: -4500px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-u3p8pb-mzNpsf { left: 0px; top: -10622px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-iBxYy-Pv6Am { left: 0px; top: -4862px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-DyVDA-r9oPif { left: -26px; top: -4774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-dZssN-D5MPn { left: 0px; top: -4780px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-LkdAo-mPlZac { left: 0px; top: -2550px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-oSWire-r9oPif { left: 0px; top: -6606px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HB1eCd-F9IAbd-OVkoRd-yaNpec { left: -20px; top: -2134px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-r9oPif { left: -26px; top: -2046px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-r9oPif-HLvlvd { left: -48px; top: -3616px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-uPjwvb-RvIlWb { left: -52px; top: -12526px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-HLvlvd { left: -40px; top: -12082px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-zMQiGf-WAutxc { left: -40px; top: -10506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-SeDgR-V7AMae { left: -62px; top: -11364px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-t5jYtc-appOce { left: -46px; top: -4374px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe-V7AMae { left: -26px; top: -12308px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DUGJie-appOce { left: 0px; top: -4984px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-aIWppb-htvI8d-r9oPif { left: -52px; top: -6538px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c { left: -40px; top: -2242px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-bOjP2c-u014N-ImhxVb-aTv5jf { left: -42px; top: -10112px; }

.HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop { left: 0px; top: -688px; }

.HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-SIsrTd { left: 0px; top: -436px; }

.HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-B1neQd-i2RYZ { left: 0px; top: -10778px; }

.HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-B1neQd-i2RYZ-SIsrTd { left: 0px; top: -6782px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nupQLb-J42Xof-zVpoTe { left: -40px; top: -1478px; }

.HB1eCd-HzV7m .HB1eCd-TIHSC-r9oPif { left: 0px; top: -2402px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TDvtud { left: -20px; top: -6856px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R { left: -14px; top: -5926px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-rymPhb-Jn51gd-r9oPif { left: 0px; top: -4754px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb-E3DyYd { left: 0px; top: -1040px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd-E3DyYd { left: -42px; top: -794px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-ZdbLkb { left: -52px; top: -7798px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-x5cW0b-E3DyYd { left: 0px; top: -12860px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-E3DyYd { left: 0px; top: -10334px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-VtOx3e-E3DyYd { left: -22px; top: -10978px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-MFS4be-E3DyYd-LSK72c { left: -61px; top: -504px; }

.HB1eCd-HzV7m .HB1eCd-DcLNVc-Xhs9z-E3DyYd { left: -42px; top: -5216px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-wUN2c-E3DyYd { left: 0px; top: -794px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-IAXTZb-E3DyYd { left: 0px; top: -9374px; }

.HB1eCd-HzV7m .HB1eCd-Yygnk-E3DyYd { left: 0px; top: -2896px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-E3DyYd { left: -20px; top: -6654px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-UlP5cd-E3DyYd { left: -26px; top: -8572px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HB1eCd-DJPBic { left: 0px; top: -10738px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-a1e4Ad-DJPBic { left: 0px; top: -1396px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RFAvhb-DJPBic { left: -60px; top: -12360px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Poonxc-eEGnhe { left: -20px; top: -1678px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Poonxc-eEGnhe-r9oPif { left: -52px; top: -4796px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nyE0bc-r9oPif { left: -46px; top: -2482px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-E3DyYd { left: -58px; top: -11900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-E3DyYd { left: -22px; top: -10736px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-E3DyYd { left: -42px; top: -7104px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-hgHJW-E3DyYd { left: -26px; top: -9420px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-OCFbXc-E3DyYd { left: 0px; top: -9694px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-z5C9Gb-E3DyYd { left: -52px; top: -10848px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xl07Ob-E3DyYd { left: -20px; top: -7512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-jNm5if-MFS4be-E3DyYd { left: -46px; top: -4334px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-OiiCO-E3DyYd { left: 0px; top: -8104px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-nUpftc-E3DyYd { left: 0px; top: -4800px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-nUpftc-MFS4be-E3DyYd { left: -40px; top: -11694px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-MFS4be-ETmUib { left: 0px; top: -2918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-E3DyYd { left: -26px; top: -5362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-KqJenf-nllRtd-E3DyYd { left: -38px; top: -6276px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-uPjwvb-ZdbLkb { left: -26px; top: -7772px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-IT5dJd-XxIAqe-E3DyYd { left: 0px; top: -3202px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-E3DyYd { left: -20px; top: -10668px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-xAa0Lb-ShBeI-E3DyYd { left: -40px; top: -5660px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Fs2VSc-r9oPif { left: 0px; top: -7772px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TNZ3Zd { left: -62px; top: -11838px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TNZ3Zd-r9oPif { left: -52px; top: -582px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec { left: 0px; top: -1698px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-jCCvxc-HNJgkc { left: -60px; top: -4650px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Bpn8Yb-E3DyYd { left: 0px; top: -11324px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif { left: 0px; top: -6520px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-UlP5cd, .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-UlP5cd { left: 0px; top: -11550px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-JbbQac-E3DyYd { left: -22px; top: -7490px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-kWbB0e-kWTbQe-E3DyYd { left: -46px; top: -3778px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-n5AaSd-E3DyYd { left: -52px; top: -10730px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rsbfue-E3DyYd { left: -46px; top: -9232px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-hxXJme-E3DyYd { left: 0px; top: -1230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ayzxhb-XPtOyb-r9oPif { left: -26px; top: -11022px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-PLDbbf-Ysl7Fe-XZYQce { left: 0px; top: -10356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-PLDbbf-SIsrTd-Ysl7Fe-XZYQce { left: 0px; top: -3382px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-DARUcf-n5AaSd-Ysl7Fe-XZYQce { left: -22px; top: -5804px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-DARUcf-n5AaSd-SIsrTd-Ysl7Fe-XZYQce { left: -26px; top: -5146px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-NGme3c-yY4Wcc-E3DyYd { left: 0px; top: -8770px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-eEDwDf-xSh02c-E3DyYd { left: 0px; top: -11000px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XPtOyb-VFQeR-E3DyYd { left: -22px; top: -8812px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-kWbB0e-kWTbQe-E3DyYd { left: 0px; top: -1778px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-ltEGzf-E3DyYd { left: 0px; top: -12022px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-RPzgNd-E3DyYd { left: 0px; top: -9446px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-i8xkGf-E3DyYd { left: 0px; top: -7624px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-fmcmS-E3DyYd { left: -58px; top: -2570px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-E3DyYd { left: 0px; top: -3616px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-E3DyYd { left: -26px; top: -6540px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-MFS4be-E3DyYd { left: -42px; top: -3512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-FMODoe-E3DyYd { left: -46px; top: -10012px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-LkdAo-E3DyYd { left: 0px; top: -1820px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-LkdAo-MFS4be-E3DyYd { left: -48px; top: -12162px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-dajHKf-E3DyYd { left: 0px; top: -4442px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-dajHKf-MFS4be-E3DyYd { left: -52px; top: -10826px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-BaYisc-E3DyYd { left: -26px; top: -9880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-BaYisc-MFS4be-E3DyYd { left: -60px; top: -1438px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-E3DyYd { left: -44px; top: -9586px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-E3DyYd { left: -20px; top: -10290px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-MFS4be-E3DyYd { left: -40px; top: -6742px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-FMODoe-E3DyYd { left: 0px; top: -1416px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-LkdAo-E3DyYd { left: -22px; top: -1348px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-LkdAo-MFS4be-E3DyYd { left: -60px; top: -1544px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-dajHKf-E3DyYd { left: -60px; top: -9184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-dajHKf-MFS4be-E3DyYd { left: 0px; top: -9586px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-BaYisc-E3DyYd { left: -44px; top: -11000px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-BaYisc-MFS4be-E3DyYd { left: 0px; top: -12184px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TDvtud-r9oPif { left: -22px; top: -9608px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-E3DyYd-EnQdTb { left: -26px; top: -7078px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-hPL1Ee-Ysl7Fe-XZYQce { left: -26px; top: -882px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-hPL1Ee-SIsrTd-Ysl7Fe-XZYQce { left: 0px; top: -10826px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-LK5yu-JeMQb { left: 0px; top: -12594px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-oXtfBe-JeMQb { left: 0px; top: -7262px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-qwU8Me-JeMQb { left: 0px; top: -11150px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-LK5yu-JeMQb { left: 0px; top: -1958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-JeMQb { left: 0px; top: -5730px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-qwU8Me-JeMQb { left: 0px; top: -8940px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-LK5yu-JeMQb { left: 0px; top: -2262px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-oXtfBe-JeMQb { left: 0px; top: -96px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-qwU8Me-JeMQb { left: 0px; top: -362px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-LK5yu-t5QKTe { left: 0px; top: -8266px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-oXtfBe-t5QKTe { left: 0px; top: -2570px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-qwU8Me-t5QKTe { left: 0px; top: -5278px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-LK5yu-t5QKTe { left: 0px; top: -736px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-t5QKTe { left: 0px; top: -6068px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-qwU8Me-t5QKTe { left: 0px; top: -12250px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-LK5yu-t5QKTe { left: 0px; top: -4192px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-oXtfBe-t5QKTe { left: -22px; top: -4442px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-qwU8Me-t5QKTe { left: -20px; top: -1172px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-LK5yu-KW5YQd-JeMQb { left: 0px; top: -6938px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-oXtfBe-KW5YQd-JeMQb { left: 0px; top: -1584px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-qwU8Me-KW5YQd-JeMQb { left: 0px; top: -3922px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-efjR6d-TzA9Ye-JeMQb { left: 0px; top: -7930px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-efjR6d-i8xkGf-JeMQb { left: 0px; top: -7698px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-aP0wEc-JeMQb { left: 0px; top: -8004px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-LK5yu-JeMQb { left: 0px; top: -5534px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-qwU8Me-JeMQb { left: 0px; top: -3704px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-s2ctBd-E3DyYd { left: -26px; top: -530px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-r9oPif { left: 0px; top: -8624px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-w9NWI-r9oPif { left: -26px; top: -10690px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-z5C9Gb { left: 0px; top: -5708px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-OCFbXc { left: 0px; top: -3996px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-tJHJj { left: -60px; top: -76px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-tJHJj-r9oPif { left: -40px; top: -9014px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-tJHJj { left: -20px; top: -7356px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-tJHJj-r9oPif { left: -52px; top: -7378px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-J9pn5c-r9oPif { left: 0px; top: -5874px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-J9pn5c-r9oPif { left: 0px; top: -12774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd-E3DyYd { left: -40px; top: -6850px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd-MFS4be-E3DyYd { left: -22px; top: -9586px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-t0O9Gd-XpSwdc { left: -42px; top: -1130px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-lxyxlb-XpSwdc { left: 0px; top: -10228px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-MFS4be-ZdbLkb { left: -52px; top: -11062px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-MFS4be-uPjwvb-ZdbLkb { left: -26px; top: -1912px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GhbEaf-xFQqWe-RvIlWb { left: -52px; top: -3228px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-ZdbLkb { left: -34px; top: -5946px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-uPjwvb-ZdbLkb { left: 0px; top: -4628px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-RvIlWb { left: 0px; top: -10072px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-uPjwvb-RvIlWb { left: 0px; top: -6336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-yqoORe-XpSwdc { left: -20px; top: -12082px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-yqoORe-RvIlWb { left: -20px; top: -4890px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-Jw1b8-uPjwvb-r9oPif { left: -22px; top: -8104px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-XPtOyb-VFQeR-XpSwdc { left: -20px; top: -2918px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-ZdbLkb { left: -20px; top: -8454px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-ZdbLkb { left: 0px; top: -1370px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nLfZJb-r9oPif { left: 0px; top: -9880px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fcEm8e-r9oPif { left: -56px; top: -5926px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-CSqGDb-yaNpec { left: 0px; top: -2336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-E3DyYd { left: -60px; top: -4292px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-CSqGDb-r9oPif { left: -26px; top: -12774px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nctj2d-yaNpec { left: -26px; top: -2376px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nctj2d-E3DyYd { left: -60px; top: -2222px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-g5XWbe-yaNpec { left: -20px; top: -8712px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-g5XWbe-r9oPif { left: 0px; top: -7818px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-KbLeYb-E3DyYd { left: -26px; top: -1034px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LUSEYe { left: 0px; top: -11900px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-LUSEYe-J9pn5c-r9oPif { left: 0px; top: -2154px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-h1U9Be { left: -62px; top: -12958px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-h1U9Be-J9pn5c-r9oPif { left: -20px; top: -816px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-HLvlvd-r9oPif { left: -22px; top: -9718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-HLvlvd-r9oPif { left: -52px; top: -9512px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-HLvlvd-i5vt6e-r9oPif { left: 0px; top: 0px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-HLvlvd-i5vt6e-r9oPif { left: -26px; top: -9828px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-mrxPge-r9oPif { left: 0px; top: -3254px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-mrxPge-r9oPif { left: 0px; top: -12334px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-mrxPge-i5vt6e-r9oPif { left: 0px; top: -1846px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-mrxPge-i5vt6e-r9oPif { left: -22px; top: -9446px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-h9d3hd-E3DyYd { left: -48px; top: -1396px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-Vkfede-ZdbLkb { left: 0px; top: -3466px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-n9oEIb-ZdbLkb { left: 0px; top: -9718px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P8wAXc-wcotoc-XzMRXd-XpSwdc { left: -52px; top: -8898px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-P8wAXc-wcotoc-XzMRXd-RvIlWb { left: 0px; top: -1518px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc-RvIlWb { left: 0px; top: -12728px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-hFsbo-XpSwdc { left: -42px; top: -3280px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-hFsbo-HLvlvd-XpSwdc { left: -20px; top: -12506px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HvfI2b-XpSwdc { left: -42px; top: -3862px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-HvfI2b-HLvlvd-XpSwdc { left: -22px; top: -794px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-uPjwvb-ZdbLkb { left: -22px; top: -11838px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-uPjwvb-RvIlWb { left: -52px; top: -6336px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-RvIlWb { left: -26px; top: -1846px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-ZdbLkb { left: 0px; top: -11716px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-XpSwdc { left: 0px; top: -12230px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c-E3DyYd { left: 0px; top: -4400px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c-r9oPif { left: 0px; top: -10446px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-FFXbQc-ZdbLkb { left: -26px; top: -8432px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc-XpSwdc { left: 0px; top: -8536px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW-XpSwdc { left: -40px; top: -4060px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ImhxVb-nMj4jb-xFQqWe-ZdbLkb { left: 0px; top: -278px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-ImhxVb-nMj4jb-MFS4be-ZdbLkb { left: -52px; top: -6584px; }

.HB1eCd-HzV7m .HB1eCd-Bz112c-DJPBic-v3pZbf-ZdbLkb { left: -20px; top: -4020px; }

.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf { background-color: white; border-top: 1px solid rgb(217, 217, 217); box-sizing: border-box; height: calc(100% - 60px); position: absolute; right: 0px; top: 60px; width: 56px; z-index: 1; }

.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf-qAWA2 { width: 0px; z-index: 1001; }

.HB1eCd-HzV7m.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf { height: calc(100% - 64px); top: 64px; }

.HB1eCd-HzV7m.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf-qAWA2 { width: 0px; }

.HB1eCd-Kk7lMc-DWWcKd-OomVLb-haAclf.HB1eCd-DWWcKd-OomVLb-haAclf-L6cTce { display: none; }

.Kk7lMc-pHHuId-b0t70b-LgbsSe.DWWcKd-OomVLb-LgbsSe { bottom: 0px; position: absolute; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-tJHJj, .Kk7lMc-pHHuId-b0t70b-xl07Ob-fmcmS { color: rgb(60, 64, 67); }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-tJHJj { font-size: 18px; font-weight: 500; line-height: 24px; padding: 6px 24px 2px; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-hgDUwe { border-top: 1px solid rgb(241, 243, 244); margin: 8px 0px; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b { border: none; cursor: pointer; height: 48px; padding: 0px; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b-sn54Q { background: rgb(241, 243, 244); }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b-Bz112c-haAclf { height: 20px; padding: 14px 16px 14px 24px; position: absolute; width: 20px; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b-OWB6Me .Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b-Bz112c { fill: rgb(218, 220, 224); }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-fmcmS { font-size: 14px; letter-spacing: 0.2px; line-height: 20px; padding: 13px 24px 11px 60px; }

.Kk7lMc-pHHuId-b0t70b-xl07Ob-ibnC6b-OWB6Me .Kk7lMc-pHHuId-b0t70b-xl07Ob-fmcmS { color: rgb(218, 220, 224); cursor: default; }

.Kk7lMc-DWWcKd-OomVLb-haAclf { background-color: white; border-left: 1px solid rgb(218, 220, 224); box-sizing: border-box; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; height: 100%; position: relative; width: 56px; }

.Kk7lMc-DWWcKd-OomVLb-Ku9FSb-haAclf { display: flex; -webkit-box-flex: 1; flex: 1 0 auto; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; margin-bottom: 56px; }

.Kk7lMc-DWWcKd-OomVLb-htvI8d-IT5dJd-haAclf { display: flex; -webkit-box-flex: 0; flex: 0 1 100%; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; padding-top: 16px; }

.Kk7lMc-DWWcKd-OomVLb-hgDUwe, .Kk7lMc-DWWcKd-OomVLb-htvI8d-IT5dJd-haAclf::before { border-top: 1px solid rgb(218, 220, 224); content: ""; display: block; -webkit-box-flex: 1; flex: 1 0 auto; margin: 0px auto; padding-bottom: 16px; width: 20px; }

.Kk7lMc-DWWcKd-OomVLb-hgDUwe { margin-top: 16px; }

.Kk7lMc-Ia7Qfc-to915.Kk7lMc-DWWcKd-OomVLb-haAclf, .Kk7lMc-Ia7Qfc-CZjX4e.Kk7lMc-DWWcKd-OomVLb-haAclf { background-color: transparent; }

.Kk7lMc-Ia7Qfc-to915.Kk7lMc-DWWcKd-OomVLb-haAclf, .Kk7lMc-Ia7Qfc-to915 .Kk7lMc-DWWcKd-OomVLb-hgDUwe, .Kk7lMc-Ia7Qfc-to915 .Kk7lMc-DWWcKd-OomVLb-htvI8d-IT5dJd-haAclf::before { border-color: rgba(255, 255, 255, 0.12); }

.Kk7lMc-Ia7Qfc-CZjX4e.Kk7lMc-DWWcKd-OomVLb-haAclf, .Kk7lMc-Ia7Qfc-CZjX4e .Kk7lMc-DWWcKd-OomVLb-hgDUwe, .Kk7lMc-Ia7Qfc-CZjX4e .Kk7lMc-DWWcKd-OomVLb-htvI8d-IT5dJd-haAclf::before { border-color: rgba(100, 121, 143, 0.12); }

.Kk7lMc-Ku9FSb-DWWcKd-OomVLb { -webkit-box-flex: 1; flex-grow: 1; height: 100px; outline: none; overflow: hidden; }

.Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge { padding: 16px 0px; }

.Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge-ojAhob { animation: 1s ease-in-out 0s infinite normal both running dotLoadingAnimation; height: 8px; background-color: rgb(117, 117, 117); border-radius: 50%; margin: 0px auto 12px; width: 8px; }

.Kk7lMc-Ia7Qfc-to915 .Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge-ojAhob { background-color: rgb(255, 255, 255); }

.Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge-ojAhob:last-child { margin-bottom: 0px; }

.Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge-ojAhob-R6PoUb { animation-delay: -0.5s; }

.Kk7lMc-DWWcKd-OomVLb-ge6pde-uDEFge-ojAhob-ibL1re { animation-delay: -0.25s; }

@-webkit-keyframes dotLoadingAnimation { 
  0%, 80%, 100% { opacity: 0.5; }
  40% { opacity: 1; }
}

@keyframes dotLoadingAnimation { 
  0%, 80%, 100% { opacity: 0.5; }
  40% { opacity: 1; }
}

.DWWcKd-OomVLb-LgbsSe { cursor: pointer; height: 56px; outline: none; pointer-events: none; position: relative; transition: all 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s; width: 56px; }

.DWWcKd-OomVLb-LgbsSe-OWB6Me { cursor: default; opacity: 0.38; }

.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .DWWcKd-OomVLb-LgbsSe-XpnDCe.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-FNFY6c .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(232, 234, 237); }

.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .DWWcKd-OomVLb-LgbsSe-FNFY6c .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(241, 243, 244); }

.Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-gk6SMd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgba(255, 255, 255, 0.24); }

.Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-FNFY6c .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-gk6SMd.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgba(255, 255, 255, 0.12); }

.DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf { background-color: transparent; background-repeat: no-repeat; background-position: center center; background-size: 20px 20px; border-radius: 50%; display: flex; -webkit-box-align: center; align-items: center; height: 40px; left: 8px; pointer-events: auto; position: absolute; top: 8px; transition: all 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s; width: 40px; }

.DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { border-radius: 50%; display: flex; height: 40px; left: 8px; position: absolute; top: 8px; transition: all 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s; width: 40px; }

.DWWcKd-OomVLb-LgbsSe-Bz112c { display: block; fill: rgb(95, 99, 104); margin: auto; transition: all 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.Kk7lMc-Ia7Qfc-to915 .DWWcKd-OomVLb-LgbsSe-Bz112c { fill: rgb(255, 255, 255); }

.DWWcKd-OomVLb-LgbsSe-zfbKYe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc.DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { animation: 3s cubic-bezier(0.05, 0.69, 0.67, 1) 0s infinite normal none running presence-scale-inner; height: 32px; width: 32px; left: 12px; top: 12px; }

.DWWcKd-OomVLb-LgbsSe-zfbKYe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc.DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { animation: 3s cubic-bezier(0.05, 0.69, 0.67, 1) 0s infinite normal none running presence-scale-outer; background-color: transparent; border-style: solid; border-width: 4px; height: 40px; width: 40px; left: 4px; top: 4px; }

.DWWcKd-OomVLb-LgbsSe-mWkOW .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc.DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { animation: 2s cubic-bezier(0.05, 0.69, 0.67, 1) 0s infinite normal none running inksplash-scale-background; }

.DWWcKd-OomVLb-LgbsSe-mWkOW .DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf { animation: 2s cubic-bezier(0.05, 0.69, 0.67, 1) 0s infinite normal none running inksplash-scale-icon; }

@-webkit-keyframes presence-scale-inner { 
  0% { opacity: 0; transform: scale(0.57); visibility: hidden; }
  15% { opacity: 0; transform: scale(0.57); visibility: visible; }
  35% { opacity: 1; transform: scale(1); }
  60% { opacity: 0; transform: scale(0.57); }
  100% { opacity: 0; transform: scale(0.57); visibility: hidden; }
}

@keyframes presence-scale-inner { 
  0% { opacity: 0; transform: scale(0.57); visibility: hidden; }
  15% { opacity: 0; transform: scale(0.57); visibility: visible; }
  35% { opacity: 1; transform: scale(1); }
  60% { opacity: 0; transform: scale(0.57); }
  100% { opacity: 0; transform: scale(0.57); visibility: hidden; }
}

@-webkit-keyframes presence-scale-outer { 
  0% { opacity: 0; transform: scale(0.75); visibility: hidden; }
  34% { opacity: 0; transform: scale(0.75); visibility: visible; }
  36% { opacity: 0.99; }
  65% { opacity: 1; }
  90% { transform: scale(1); }
  100% { opacity: 0; transform: scale(1); visibility: hidden; }
}

@keyframes presence-scale-outer { 
  0% { opacity: 0; transform: scale(0.75); visibility: hidden; }
  34% { opacity: 0; transform: scale(0.75); visibility: visible; }
  36% { opacity: 0.99; }
  65% { opacity: 1; }
  90% { transform: scale(1); }
  100% { opacity: 0; transform: scale(1); visibility: hidden; }
}

@-webkit-keyframes inksplash-scale-background { 
  0% { opacity: 0; transform: scale(0); }
  35% { opacity: 0; transform: scale(0.4); }
  50% { opacity: 1; }
  80% { transform: scale(2.05); }
  100% { opacity: 0; transform: scale(0); }
}

@keyframes inksplash-scale-background { 
  0% { opacity: 0; transform: scale(0); }
  35% { opacity: 0; transform: scale(0.4); }
  50% { opacity: 1; }
  80% { transform: scale(2.05); }
  100% { opacity: 0; transform: scale(0); }
}

@-webkit-keyframes inksplash-scale-icon { 
  0% { transform: scale(1); }
  20% { transform: scale(1); }
  30% { transform: scale(1.1); }
  40% { transform: scale(1); }
  100% { transform: scale(1); }
}

@keyframes inksplash-scale-icon { 
  0% { transform: scale(1); }
  20% { transform: scale(1); }
  30% { transform: scale(1.1); }
  40% { transform: scale(1); }
  100% { transform: scale(1); }
}

.DWWcKd-OomVLb-xl07Ob { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.2); border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; min-width: 180px; outline: none; overflow-y: auto; padding: 8px 0px; position: absolute; z-index: 1202; }

.Kk7lMc-QWPxkf-LgbsSe-haAclf { bottom: 0px; display: flex; height: 56px; overflow: hidden; pointer-events: none; position: absolute; right: 0px; width: 56px; }

.Kk7lMc-QWPxkf-LgbsSe-haAclf.Kk7lMc-QWPxkf-LgbsSe-haAclf-uQVisb { margin-bottom: 24px; }

.Kk7lMc-QWPxkf-LgbsSe { bottom: 0px; }

.Kk7lMc-QWPxkf-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf, .Kk7lMc-QWPxkf-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { border-radius: calc(58px); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(255, 255, 255); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(241, 243, 244); }

.Kk7lMc-Ia7Qfc-to915 .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(89, 89, 89); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc, .Kk7lMc-Ia7Qfc-CZjX4e .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { background-color: rgb(232, 234, 237); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie { right: -24px; }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf { border-bottom-right-radius: 0px; border-top-right-radius: 0px; height: 20px; left: 0px; margin: 8px 0px 8px 8px; padding: 10px 0px 10px 10px; top: 0px; width: calc(58px); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { border-bottom-right-radius: 0px; border-top-right-radius: 0px; height: 20px; left: 0px; margin: 8px 0px 8px 8px; padding: 10px 0px 10px 10px; top: 0px; width: calc(58px); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 1px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-ZmdkE { right: 0px; }

.Kk7lMc-QWPxkf-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c { left: 10px; position: absolute; top: 10px; }

html[dir="rtl"] .Kk7lMc-QWPxkf-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c, body[dir="rtl"] .Kk7lMc-QWPxkf-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c { transform: rotate(180deg); }

.Kk7lMc-Ia7Qfc-to915 .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf, .Kk7lMc-Ia7Qfc-to915 .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-haAclf { background-color: rgb(65, 65, 65); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c { margin-left: -6px; transform: rotate(180deg); }

.Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c { margin-left: 0px; }

html[dir="rtl"] .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c, body[dir="rtl"] .Kk7lMc-QWPxkf-LgbsSe.DWWcKd-OomVLb-LgbsSe-barxie .DWWcKd-OomVLb-LgbsSe-Bz112c { transform: rotate(0deg); }

.VL4Fef-GIHV4-bnBfGc { background-color: white; background-repeat: no-repeat; border: transparent; border-radius: 8px; box-sizing: border-box; color: rgb(102, 102, 102); height: 56px; outline: none; padding: 0px 10px; pointer-events: none; position: fixed; z-index: 999; }

.VL4Fef-GIHV4-bnBfGc.VL4Fef-GIHV4-bnBfGc-LJTIlf-rTEl { background-position: 20px center; background-size: 24px 24px; height: 56px; width: 200px; }

.VL4Fef-GIHV4-bnBfGc.VL4Fef-GIHV4-bnBfGc-HiaYvf-rTEl { background-position: center center; background-size: 100%; height: 120px; width: 120px; }

.VL4Fef-GIHV4-bnBfGc.VL4Fef-GIHV4-bnBfGc-HiaYvf-rTEl.VL4Fef-GIHV4-bnBfGc-HiaYvf-bmhONe { height: 156px; }

.VL4Fef-GIHV4-bnBfGc-fmcmS-i8xkGf { box-sizing: border-box; display: table-cell; padding-left: 48px; max-width: 200px; vertical-align: middle; }

.VL4Fef-GIHV4-bnBfGc-fmcmS-i8xkGf .VL4Fef-GIHV4-bnBfGc-r4nke { font-size: 1.1em; }

.VL4Fef-GIHV4-bnBfGc-fmcmS-i8xkGf .VL4Fef-GIHV4-bnBfGc-fmcmS { opacity: 0.75; padding-top: 2px; }

.VL4Fef-GIHV4-bnBfGc-HiaYvf-rTEl .VL4Fef-GIHV4-bnBfGc-fmcmS { background-color: rgba(32, 33, 36, 0.71); border-radius: 0px 0px 8px 8px; bottom: 0px; color: white; height: 36px; left: 0px; padding: 8px 10px; position: absolute; width: 100%; }

.VL4Fef-GIHV4-bnBfGc .VL4Fef-GIHV4-bnBfGc-r4nke, .VL4Fef-GIHV4-bnBfGc .VL4Fef-GIHV4-bnBfGc-fmcmS { box-sizing: border-box; margin: 0px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.VL4Fef-GIHV4-bnBfGc .VL4Fef-GIHV4-bnBfGc-NnAfwf-VCkuzd { background-color: rgb(32, 33, 36); border-radius: 20px; box-sizing: border-box; color: white; font-size: 16px; height: 40px; max-width: 75%; min-width: 40px; overflow: hidden; padding: 9px 8px; position: absolute; right: -15px; text-align: center; text-overflow: ellipsis; top: -15px; }

.UPJOje-vYU7ve { height: inherit; position: relative; width: 100%; }

.UPJOje-bN97Pc { height: 100%; left: 0px; position: absolute; top: 0px; width: 100%; z-index: 0; }

.ONKrsd-jrnDlb-ho7Xm-VPIWce::after { content: ""; background-color: rgb(219, 68, 55); border-radius: 50%; height: 8px; position: absolute; right: 17px; top: 17px; width: 8px; }

.Kk7lMc-Ku9FSb-DWWcKd-OomVLb .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgb(232, 240, 254); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-v3pZbf .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgba(66, 133, 244, 0.24); }

.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgb(230, 244, 234); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgba(52, 168, 83, 0.24); }

.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgb(254, 247, 224); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgba(251, 188, 4, 0.24); }

.Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-n0tgWb { border-color: rgba(255, 255, 255, 0.24); }

.Kk7lMc-Ku9FSb-DWWcKd-OomVLb .DWWcKd-OomVLb-LgbsSe-mWkOW .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ku9FSb-DWWcKd-OomVLb .DWWcKd-OomVLb-LgbsSe-zfbKYe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ku9FSb-DWWcKd-OomVLb .DWWcKd-OomVLb-LgbsSe-gk6SMd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-v3pZbf.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(232, 240, 254); }

.DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-v3pZbf.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(210, 227, 252); }

.Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-mWkOW.ONKrsd-jrnDlb-v3pZbf .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-zfbKYe.ONKrsd-jrnDlb-v3pZbf .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-v3pZbf .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-v3pZbf.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(66, 133, 244, 0.24); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-v3pZbf.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-v3pZbf.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(66, 133, 244, 0.12); }

.DWWcKd-OomVLb-LgbsSe-mWkOW.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-zfbKYe.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-nllRtd.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(230, 244, 234); }

.DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-nllRtd.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(206, 234, 214); }

.Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-mWkOW.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-zfbKYe.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-nllRtd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-nllRtd.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(52, 168, 83, 0.24); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-nllRtd.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-nllRtd.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(52, 168, 83, 0.12); }

.DWWcKd-OomVLb-LgbsSe-mWkOW.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-zfbKYe.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-gS7Ybc.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(254, 247, 224); }

.DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-gS7Ybc.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgb(254, 239, 195); }

.Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-mWkOW.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-zfbKYe.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-gS7Ybc .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .DWWcKd-OomVLb-LgbsSe-gk6SMd.ONKrsd-jrnDlb-gS7Ybc.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(251, 188, 4, 0.24); }

.Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-gS7Ybc.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-CZjX4e .ONKrsd-jrnDlb-gS7Ybc.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(251, 188, 4, 0.12); }

.Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-mWkOW .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-zfbKYe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-gk6SMd .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-gk6SMd.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(255, 255, 255, 0.24); }

.Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-ZmdkE .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb, .Kk7lMc-Ia7Qfc-to915 .ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-XpnDCe .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc-SmKAyb { background-color: rgba(255, 255, 255, 0.12); }

.ONKrsd-jrnDlb-Bz112c-gvZm2b-uDEFge { background-color: rgb(215, 4, 251); border-radius: 3px 0px 0px 3px; display: none; height: 40px; position: absolute; right: 1px; top: 8px; width: 3px; }

.ONKrsd-jrnDlb-LgbsSe.DWWcKd-OomVLb-LgbsSe-gk6SMd .ONKrsd-jrnDlb-Bz112c-gvZm2b-uDEFge { display: inherit; }

.ONKrsd-jrnDlb-v3pZbf .ONKrsd-jrnDlb-Bz112c-gvZm2b-uDEFge { background-color: rgb(66, 133, 244); }

.ONKrsd-jrnDlb-nllRtd .ONKrsd-jrnDlb-Bz112c-gvZm2b-uDEFge { background-color: rgb(52, 168, 83); }

.ONKrsd-jrnDlb-gS7Ybc .ONKrsd-jrnDlb-Bz112c-gvZm2b-uDEFge { background-color: rgb(251, 188, 4); }

.Kk7lMc-Ia7Qfc-to915 .Kk7lMc-RPzgNd-xl07Ob-LgbsSe:not(.DWWcKd-OomVLb-LgbsSe-ZmdkE) .DWWcKd-OomVLb-LgbsSe-Bz112c-AHe6Kc { opacity: 0.7; }

.Kk7lMc-ae3xF-tJHJj { -webkit-box-align: center; align-items: center; background-color: rgb(255, 255, 255); border-bottom: 1px solid rgb(241, 243, 244); box-sizing: border-box; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: row; -webkit-font-smoothing: antialiased; height: 64px; padding: 0px 10px; position: relative; z-index: 1; }

.Kk7lMc-ae3xF-tJHJj-PQbLGe { margin-left: 10px; margin-right: 10px; }

.Kk7lMc-ae3xF-r4nke-haAclf { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex-grow: 1; -webkit-box-pack: center; justify-content: center; width: 1px; }

.Kk7lMc-ae3xF-r4nke-PQbLGe { margin: 0px; }

.Kk7lMc-ae3xF-r4nke-fmcmS, .Kk7lMc-ae3xF-VdSJob-fmcmS, .Kk7lMc-ae3xF-VdSJob-fmcmS .VIpgJd-xl07Ob-LgbsSe-cHYyed { overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.Kk7lMc-ae3xF-r4nke-fmcmS, .Kk7lMc-ae3xF-VdSJob-fmcmS { outline: none; }

.Kk7lMc-ae3xF-r4nke-fmcmS.Kk7lMc-ae3xF-r4nke-zfdrlf { font-size: 22px; }

.Kk7lMc-ae3xF-tJHJj-CZjX4e-AHe6Kc .Kk7lMc-ae3xF-r4nke-zfdrlf { color: rgba(0, 0, 0, 0.54); }

.Kk7lMc-ae3xF-tJHJj-to915-AHe6Kc .Kk7lMc-ae3xF-r4nke-zfdrlf { color: rgb(255, 255, 255); }

.Kk7lMc-ae3xF-r4nke-fmcmS.Kk7lMc-ae3xF-r4nke-purZT { color: rgb(95, 99, 104); font-size: 10px; font-weight: 500; letter-spacing: 1.5px; text-transform: uppercase; }

.Kk7lMc-ae3xF-r4nke-fmcmS.Kk7lMc-ae3xF-r4nke-purZT.Kk7lMc-ae3xF-KQ1Bvd { left: 56px; }

.Kk7lMc-ae3xF-j4gsHd-haAclf { font-size: 0px; }

.Kk7lMc-ae3xF-VdSJob-fmcmS { color: rgb(60, 64, 67); font-size: 16px; font-weight: 500; line-height: 20px; }

.Kk7lMc-ae3xF-VdSJob-fmcmS.VIpgJd-xl07Ob-LgbsSe-FNFY6c { background-color: rgb(241, 243, 244); }

.Kk7lMc-ae3xF-VdSJob-LgbsSe { padding: 0px 2px 0px 4px; }

.Kk7lMc-ae3xF-VdSJob-LgbsSe .Kk7lMc-ae3xF-VdSJob-fmcmS, .Kk7lMc-ae3xF-VdSJob-fmcmS .VIpgJd-xl07Ob-LgbsSe-cHYyed { padding: 0px; }

.Kk7lMc-ae3xF-VdSJob-F75qrd-m9bMae { color: rgb(26, 115, 232); }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe { background: none; border-radius: 3px; border-width: 0px; box-sizing: border-box; cursor: pointer; display: inline-block; margin-left: -4px; max-width: 100%; outline: none; padding: 0px 2px 0px 4px; }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe.Kk7lMc-ae3xF-j4gsHd-LgbsSe-ZmdkE { background-color: rgb(241, 243, 244); }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe.Kk7lMc-ae3xF-j4gsHd-LgbsSe-XpnDCe, .Kk7lMc-ae3xF-j4gsHd-LgbsSe.Kk7lMc-ae3xF-j4gsHd-LgbsSe-FNFY6c { background-color: rgb(232, 234, 237); }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe.Kk7lMc-ae3xF-j4gsHd-LgbsSe-OWB6Me { opacity: 0.38; }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe .Kk7lMc-ae3xF-j4gsHd-LgbsSe-n0tgWb-Q4BLdf { display: flex; justify-content: flex-start; }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe .Kk7lMc-ae3xF-j4gsHd-LgbsSe-SmKAyb-Q4BLdf { display: block; flex-shrink: 1; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.Kk7lMc-ae3xF-j4gsHd-LgbsSe-n0tgWb-Q4BLdf::after { content: ""; display: block; background: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0naHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmcnIHdpZHRoPScyNHB4JyBoZWlnaHQ9JzI0cHgnIHZpZXdCb3g9JzAgMCAyNCAyNCcgZmlsbD0nIzVmNjM2OCc+PHBhdGggZD0nTTcgMTBsNSA1IDUtNXonPjwvcGF0aD48cGF0aCBkPSdNMCAwaDI0djI0SDB6JyBmaWxsPSdub25lJz48L3BhdGg+PC9zdmc+") center center no-repeat; flex-shrink: 0; height: 20px; margin: 0px 0px 0px 4px; padding: 0px; width: 20px; }

.Kk7lMc-ae3xF-tJHJj-c6xFrd { display: flex; height: 24px; justify-content: flex-end; position: absolute; right: 8px; top: 18px; }

.Kk7lMc-ae3xF-tJHJj-LgbsSe { background: center center / 20px 20px no-repeat; cursor: pointer; height: 24px; width: 24px; }

.Kk7lMc-ae3xF-tJHJj-CZjX4e-AHe6Kc .Kk7lMc-ae3xF-tJHJj-OAU7Vd-Bz112c { fill: rgb(0, 0, 0); opacity: 0.54; }

.Kk7lMc-ae3xF-tJHJj-to915-AHe6Kc .Kk7lMc-ae3xF-tJHJj-OAU7Vd-Bz112c { fill: rgb(255, 255, 255); }

html[dir="rtl"] .Kk7lMc-ae3xF-a4fUwd-LgbsSe, body[dir="rtl"] .Kk7lMc-ae3xF-a4fUwd-LgbsSe, html[dir="rtl"] .Kk7lMc-ae3xF-FwpN6e-d5JObf-LgbsSe, body[dir="rtl"] .Kk7lMc-ae3xF-FwpN6e-d5JObf-LgbsSe { transform: scaleX(-1); }

.Kk7lMc-ae3xF-tJHJj-LgbsSe.Kk7lMc-ae3xF-r4nke-PQbLGe { margin: 0px; }

.Kk7lMc-ae3xF-tJHJj-LgbsSe:hover { opacity: 0.87; }

.Kk7lMc-ae3xF-VdSJob-LgbsSe[aria-disabled="true"], .Kk7lMc-ae3xF-tJHJj-LgbsSe[aria-disabled="true"] { cursor: not-allowed; opacity: 0.38; }

.Kk7lMc-ae3xF-a4fUwd-LgbsSe { margin-right: 2px; }

.VIpgJd-xl07Ob.Kk7lMc-ae3xF-DaY83b-hgHJW-xl07Ob { background: rgb(255, 255, 255); border-width: 0px; border-radius: 0px 0px 8px 8px; box-shadow: rgba(0, 0, 0, 0.12) 0px -3px 6px -3px, rgba(0, 0, 0, 0.14) 0px 4px 8px -2px; box-sizing: border-box; max-height: 400px; overflow: hidden auto; padding-bottom: 8px; position: absolute; width: 100%; z-index: 999; }

.VIpgJd-j7LFlb.Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd { border: none; height: 40px; padding: 0px; width: 300px; }

.VIpgJd-j7LFlb-sn54Q.Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd { background: rgb(241, 243, 244); }

.VIpgJd-xl07Ob.Kk7lMc-ae3xF-DaY83b-hgHJW-xl07Ob .VIpgJd-gqMrKb { border-top: 1px solid rgba(32, 33, 36, 0.06); margin: 8px 0px; padding: 0px; }

.Kk7lMc-ae3xF-DaY83b-hgHJW-g6cJHd { display: none; height: 20px; padding: 10px 16px; position: absolute; right: 0px; width: 20px; }

.VIpgJd-wQNmvb-gk6SMd .Kk7lMc-ae3xF-DaY83b-hgHJW-g6cJHd { display: block; }

.Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd.VIpgJd-wQNmvb-gk6SMd { background-image: none; }

.Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd .VIpgJd-j7LFlb-MPu53c, .Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd.VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-MPu53c { display: none; }

.Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd-fmcmS { box-sizing: border-box; font-size: 14px; color: rgb(32, 33, 36); padding: 10px 20px; letter-spacing: 0.2px; line-height: 20px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; width: 300px; }

.VIpgJd-wQNmvb-gk6SMd .Kk7lMc-ae3xF-DaY83b-hgHJW-x3Eknd-fmcmS { padding-right: 60px; }

.Kk7lMc-ae3xF-bN97Pc-LYNcwc { background-color: white; box-sizing: border-box; height: 100%; left: 0px; padding-top: 64px; position: absolute; top: 0px; width: 100%; }

.Kk7lMc-tJHJj-bEDTcc-L5Fo6c .Kk7lMc-ae3xF-Ku9FSb { padding-top: 0px; }

.Kk7lMc-ae3xF-ge6pde { overflow: hidden; position: absolute; text-align: center; }

.Kk7lMc-ae3xF-PrY1nf, .Kk7lMc-ae3xF-zozyIf-gcuqQc, .Kk7lMc-ae3xF-XrLSYd-m9bMae, .Kk7lMc-ae3xF-lJi4pf { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; text-align: center; }

.Kk7lMc-ae3xF-PrY1nf-ij8cu, .Kk7lMc-ae3xF-PrY1nf-r4nke, .Kk7lMc-ae3xF-lJi4pf-ij8cu, .Kk7lMc-ae3xF-lJi4pf-r4nke { color: rgb(95, 99, 104); margin: 0px 70px; }

.Kk7lMc-ae3xF-PrY1nf-ij8cu, .Kk7lMc-ae3xF-lJi4pf-ij8cu { font-size: 12px; line-height: 16px; }

.Kk7lMc-ae3xF-PrY1nf-r4nke, .Kk7lMc-ae3xF-lJi4pf-r4nke { font-size: 16px; font-weight: 500; margin-bottom: 2px; margin-top: 34px; }

.Kk7lMc-ae3xF-zozyIf-gcuqQc-Ne3sFf, .Kk7lMc-ae3xF-XrLSYd-m9bMae-Ne3sFf { margin: 10px; max-width: calc(100% - 20px); }

.Kk7lMc-ae3xF-XrLSYd-m9bMae-dTKROe { color: rgb(26, 115, 232); cursor: pointer; text-transform: uppercase; }

.Kk7lMc-ae3xF-XrLSYd-m9bMae-TZk80d-Jwxghc { margin-top: 40px; }

.Kk7lMc-ae3xF-L5Fo6c { border: 0px; height: 100%; width: 100%; }

.Kk7lMc-ae3xF-G0jgYd-haAclf { -webkit-box-align: center; align-items: center; background-color: rgb(255, 255, 255); box-sizing: border-box; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: row; height: 100%; left: 0px; padding: 0px 10px; position: absolute; top: 0px; width: 100%; }

.Kk7lMc-ae3xF-G0jgYd-Bz112c, .Kk7lMc-ae3xF-G0jgYd-TvD9Pc { margin-left: 10px; margin-right: 10px; }

.Kk7lMc-ae3xF-G0jgYd-YPqjbf { background-color: transparent; border: none; color: rgb(95, 99, 104); -webkit-box-flex: 1; flex-grow: 1; font-size: 16px; line-height: 24px; outline: none; width: 100px; }

.Kk7lMc-ae3xF-G0jgYd-YPqjbf::placeholder { color: rgb(189, 193, 198); }

.Kk7lMc-ae3xF-G0jgYd-YPqjbf::-webkit-input-placeholder { color: rgb(189, 193, 198); }

.Kk7lMc-DWWcKd-OomVLb-haAclf .tk3N6e-VCkuzd { padding: 16px; border-radius: 8px; border-color: rgb(232, 234, 237); border-width: 1px; box-shadow: rgba(60, 64, 67, 0.3) 0px 2px 6px; }

.Kk7lMc-DWWcKd-OomVLb-haAclf .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc { border-left-color: rgb(232, 234, 237); border-right-color: rgb(232, 234, 237); }

.DWWcKd-OomVLb-b3rLgd-VCkuzd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-tJHJj { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: row; height: 32px; width: 200px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-HiaYvf-haAclf { width: 32px; border-radius: 50%; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-HiaYvf-haAclf .DWWcKd-OomVLb-b3rLgd-VCkuzd-HiaYvf { width: 32px; height: 32px; border-radius: 50%; margin-right: 8px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-fmcmS { height: 31.5px; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; margin-left: 8px; margin-bottom: 8px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-fmcmS:focus { outline: none; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-r4nke-fmcmS { height: 14px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; color: rgb(95, 99, 104); }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-qJTHM-fmcmS { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; color: rgb(60, 64, 67); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-yePe5c { margin-top: 9px; height: 32px; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: row; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-yePe5c .tk3N6e-LgbsSe { text-align: center; font-weight: 500; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding-left: 8px; padding-right: 16px; margin: 0px; height: 30px; line-height: 30px; color: rgb(255, 255, 255); max-width: 300px; font-size: 14px; border-radius: 15px; -webkit-box-align: center; align-items: center; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-yePe5c .DWWcKd-OomVLb-b3rLgd-VCkuzd-LgbsSe-Bz112c { width: 16px; height: 16px; padding-right: 8px; padding-top: 6px; padding-bottom: 7px; vertical-align: middle; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-yePe5c .DWWcKd-OomVLb-b3rLgd-VCkuzd-DbgRPb { width: 8px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-F75qrd-wcotoc-JIbuQc-LgbsSe { background-color: rgb(24, 128, 56); }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-F75qrd-wcotoc-JIbuQc-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(42, 137, 71); box-shadow: rgba(24, 128, 56, 0.15) 0px 1px 3px 1px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-F75qrd-wcotoc-JIbuQc-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background-color: rgb(79, 158, 103); box-shadow: rgba(24, 128, 56, 0.15) 0px 1px 3px 1px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-F75qrd-wcotoc-JIbuQc-LgbsSe.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(98, 168, 119); box-shadow: rgba(24, 128, 56, 0.15) 0px 1px 3px 1px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-IYtByb-LgbsSe { background-color: rgb(217, 48, 37); }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-IYtByb-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(211, 68, 59); box-shadow: rgba(217, 48, 37, 0.15) 0px 1px 3px 1px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-IYtByb-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background-color: rgb(224, 108, 100); box-shadow: rgba(217, 48, 37, 0.15) 0px 1px 3px 1px; }

.DWWcKd-OomVLb-b3rLgd-VCkuzd .DWWcKd-OomVLb-b3rLgd-VCkuzd-IYtByb-LgbsSe.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(232, 138, 132); box-shadow: rgba(217, 48, 37, 0.15) 0px 1px 3px 1px; }

.Kk7lMc-RPzgNd-xl07Ob-ibnC6b { -webkit-box-align: center; align-items: center; cursor: pointer; display: flex; padding: 8px; }

.Kk7lMc-RPzgNd-xl07Ob-ibnC6b-sn54Q { background-color: rgb(241, 243, 244); }

.Kk7lMc-RPzgNd-xl07Ob-ibnC6b-Bz112c { background: center center / 20px 20px no-repeat transparent; border-radius: 50%; height: 40px; width: 40px; }

.Kk7lMc-RPzgNd-xl07Ob-ibnC6b-bN97Pc { padding: 0px 6px; white-space: nowrap; }

.Kk7lMc-RPzgNd-xl07Ob-ibnC6b-OWB6Me { cursor: default; opacity: 0.38; }

.Kk7lMc-FbH7jb-rcuQ6b .UPJOje-bN97Pc { animation: 333ms ease 0s 1 normal both paused companion-server-render-guest-content-fadeout; }

.Kk7lMc-FbH7jb-rcuQ6b .Kk7lMc-ae3xF-jgixuf-uMX1Ee-kWbB0e-jgixuf-hxXJme { display: none; }

.Kk7lMc-FbH7jb-rcuQ6b .Kk7lMc-ae3xF-jgixuf-uMX1Ee-DWWcKd-l4eHX { animation: 0s ease 0s 1 normal none running none; }

.Kk7lMc-FbH7jb-rcuQ6b .Kk7lMc-ae3xF-jgixuf-uMX1Ee-jH4Ejd { display: none; }

@-webkit-keyframes companion-server-render-guest-content-fadeout { 
  0% { opacity: 0.38; }
  100% { opacity: 0; }
}

@keyframes companion-server-render-guest-content-fadeout { 
  0% { opacity: 0.38; }
  100% { opacity: 0; }
}

.Kk7lMc-ae3xF { background-color: white; box-sizing: border-box; height: 100%; width: 300px; }

.Kk7lMc-ae3xF:not(.Kk7lMc-FbH7jb-rcuQ6b) { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; }

.Kk7lMc-ae3xF-WdRn2-bN97Pc-haAclf, .Kk7lMc-ae3xF-Ku9FSb-bN97Pc-haAclf, .Kk7lMc-ae3xF-MVH0Ye-bN97Pc-haAclf { height: 100%; }

.Kk7lMc-ae3xF.Kk7lMc-ae3xF-bF1uUb-bN97Pc { border: 0px; box-shadow: rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px, rgba(0, 0, 0, 0.2) 0px 2px 4px -1px; opacity: 1; }

.Kk7lMc-ae3xF-DWWcKd-OomVLb { bottom: 0px; left: 0px; position: absolute; }

.Kk7lMc-ae3xF-Ku9FSb-haAclf { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; height: 100%; }

.Kk7lMc-ae3xF-jgixuf-uMX1Ee-haAclf { height: 680px; margin-left: 50%; position: relative; top: calc(50% - 404px); transform: translateX(-50%); width: 680px; }

html[dir="rtl"] .Kk7lMc-ae3xF-jgixuf-uMX1Ee-haAclf, body[dir="rtl"] .Kk7lMc-ae3xF-jgixuf-uMX1Ee-haAclf { transform: translateX(50%); }

.Kk7lMc-ae3xF-jgixuf-uMX1Ee-kWbB0e-jgixuf-hxXJme { animation: 1s cubic-bezier(0.08, 0.8, 0.67, 1) 400ms 1 normal both running ink-splash-opacity, 1s cubic-bezier(0.05, 0.69, 0.67, 1) 400ms 1 normal both running ink-splash-scale; border-radius: 50%; height: 100%; width: 100%; }

@-webkit-keyframes ink-splash-opacity { 
  0% { opacity: 1; }
  100% { opacity: 0; }
}

@keyframes ink-splash-opacity { 
  0% { opacity: 1; }
  100% { opacity: 0; }
}

@-webkit-keyframes ink-splash-scale { 
  0% { transform: scale(0); }
  100% { transform: scale(1); }
}

@keyframes ink-splash-scale { 
  0% { transform: scale(0); }
  100% { transform: scale(1); }
}

.Kk7lMc-ae3xF-jgixuf-uMX1Ee-DWWcKd-l4eHX { animation: 330ms cubic-bezier(0.05, 0.62, 0.51, 1.26) 333ms 1 normal backwards running app-logo-scale, 170ms cubic-bezier(0.29, 0, 0.73, 1) 667ms 1 normal forwards running app-logo-scale-bounce; background-position: center center; background-repeat: no-repeat; background-size: 128px 128px; inset: 0px; height: 128px; margin: auto; position: absolute; width: 128px; }

@-webkit-keyframes app-logo-scale { 
  0% { transform: scale(0); }
  100% { transform: scale(1); }
}

@keyframes app-logo-scale { 
  0% { transform: scale(0); }
  100% { transform: scale(1); }
}

@-webkit-keyframes app-logo-scale-bounce { 
  0%, 100% { transform: scale(1); }
  20% { transform: scale(0.95); }
}

@keyframes app-logo-scale-bounce { 
  0%, 100% { transform: scale(1); }
  20% { transform: scale(0.95); }
}

.Kk7lMc-ae3xF-jgixuf-uMX1Ee-jH4Ejd { animation: 330ms linear 1s 1 normal both running beachball-opacity; inset: 190px 0px 0px; height: 20px; margin: auto; position: absolute; width: 20px; }

@-webkit-keyframes beachball-opacity { 
  0% { opacity: 0; }
  100% { opacity: 1; }
}

@keyframes beachball-opacity { 
  0% { opacity: 0; }
  100% { opacity: 1; }
}

.Kk7lMc-suEOdc { background-color: rgba(60, 64, 67, 0.9); border-radius: 4px; color: rgb(255, 255, 255); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 500; -webkit-font-smoothing: antialiased; letter-spacing: 0.3px; line-height: 16px; padding: 4px 8px; white-space: nowrap; z-index: 9999; }

.HB1eCd-Kk7lMc-PvRhvb { box-shadow: rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px, rgba(0, 0, 0, 0.2) 0px 2px 4px -1px; height: 100%; outline: none; overflow: hidden; position: absolute; right: 0px; top: 0px; width: 300px; z-index: 901; }

.HB1eCd-Qrtp3c-yBi6gb { -webkit-user-drag: none; user-select: none; }

#docs-chrome { background: white; outline: none; }

#docs-chrome.HB1eCd-R1gDOc-NMrWyd { border-bottom: 1px solid rgb(217, 217, 217); min-height: 56px; }

#docs-header { position: relative; flex: 1 1 auto; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb { height: 49px; }

#docs-header.HB1eCd-aSVJYc-x5AlNc { max-height: 31px; }

#docs-header-container, #docs-banner-container { display: flex; justify-content: flex-end; }

#docs-banners { overflow: hidden; position: relative; flex: 1 1 auto; }

#docs-account-level-banner { display: flex; white-space: nowrap; width: 100%; }

#docs-file-level-banner { display: flex; flex-direction: column; white-space: nowrap; width: 100%; }

.HB1eCd-Vkfede-NBtyUd-PvRhvb-LwH6nd { flex: 0 0 0px; }

.HB1eCd-Vkfede-NBtyUd-PvRhvb-LwH6nd.PBWx0c { flex-basis: 300px; }

.HB1eCd-PvRhvb-tJHJj-fmcmS { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; left: 20px; position: absolute; font-size: 14px; }

.HB1eCd-PvRhvb-gGtCd { overflow: hidden; }

#docs-bars { position: relative; }

#docs-titlebar-container { margin-left: 40px; position: relative; }

#docs-branding-container { height: 60px; margin-top: 26px; position: absolute; width: 40px; z-index: 1; }

#docs-branding-container a { display: inline-block; height: 60px; width: 40px; }

.HB1eCd-aSVJYc-x5AlNc #docs-branding-container { margin-top: 0px; }

.HB1eCd-HzV7m #docs-branding-container #docs-branding-ehb { cursor: pointer; height: 0px; left: 8px; margin: unset; padding: unset; position: absolute; transform: rotate(-45deg) translateX(-14px); top: 20px; width: unset; z-index: 1; }

[dir="rtl"] .HB1eCd-HzV7m #docs-branding-container #docs-branding-ehb { transform: rotate(45deg) translateX(14px); }

#docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-fmcmS { color: rgb(255, 255, 255); font-weight: 500; left: 8px; position: absolute; top: 5px; z-index: 1; }

#docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-bRIwWb { border-radius: 2px; height: 22px; position: absolute; transform: perspective(29px) rotateX(49deg); width: 50px; }

.HB1eCd-n7vHCb-arrpzb #docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-fmcmS { color: rgb(0, 0, 0); }

.HB1eCd-n7vHCb-arrpzb #docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-bRIwWb { background: rgb(255, 149, 0); }

.HB1eCd-n7vHCb-TftRv #docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-bRIwWb { background: rgb(0, 102, 218); }

.HB1eCd-n7vHCb-G1jlMc #docs-branding-ehb .HB1eCd-n7vHCb-NoGbpc-bRIwWb { background: rgb(0, 131, 45); }

#docs-titlebar { clear: both; font-size: 18px; height: 24px; padding: 7px 0px 0px; width: 100%; }

.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar { font-size: 16px; }

#docs-header.HB1eCd-aSVJYc-x5AlNc #docs-titlebar { height: 24px; padding-top: 0px; }

#docs-header.HB1eCd-aSVJYc-x5AlNc #docs-titlebar-container { top: -21px; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-container { height: 100%; }

#docs-header.HB1eCd-aSVJYc-x5AlNc .HB1eCd-NezmJd-c6xFrd { top: 19px; }

.HB1eCd-rcyUVe { border-radius: 6px; border: 1px solid rgb(136, 0, 0); color: rgb(136, 0, 0); float: left; font-size: 11px; margin-right: 8px; padding: 0px 5px; text-align: center; white-space: nowrap; }

#docs-drive-logo { height: 60px; position: absolute; width: 40px; opacity: 0; transition: all 125ms linear 0s; }

#docs-branding-logo { height: 60px; position: absolute; width: 40px; transition: all 125ms linear 0s; }

#docs-branding-container.HB1eCd-n7vHCb-zTETae { background-color: rgb(209, 209, 209); }

#docs-branding-container.HB1eCd-n7vHCb-TftRv { background-color: rgb(66, 133, 244); }

#docs-branding-container.HB1eCd-n7vHCb-G1jlMc { background-color: rgb(15, 157, 88); }

#docs-branding-container.HB1eCd-n7vHCb-arrpzb { background-color: rgb(244, 180, 0); }

#docs-branding-container.HB1eCd-n7vHCb-QymXn { background-color: rgb(219, 68, 55); }

#docs-branding-container.HB1eCd-n7vHCb-t02dhe { background-color: rgb(103, 58, 183); }

#docs-branding-container.HB1eCd-n7vHCb-jdTLZc { background-color: rgb(66, 133, 244); }

#docs-branding-container:not(.HB1eCd-n7vHCb-OQ09Xb-RCfa3e-OWB6Me):hover #docs-drive-logo { opacity: 1; }

#docs-branding-container:not(.HB1eCd-n7vHCb-OQ09Xb-RCfa3e-OWB6Me):hover #docs-branding-logo { opacity: 0; }

#docs-branding-container.HB1eCd-n7vHCb-zTETae:hover #docs-drive-logo { opacity: 0; }

#docs-branding-container.HB1eCd-n7vHCb-zTETae:hover #docs-branding-logo { opacity: 1; }

.HB1eCd-PLEiK { text-align: center; }

.HB1eCd-PLEiK-SmKAyb { border-radius: 3px; font-size: 13px; font-weight: 500; margin: 0px auto 5px; padding: 5px 7px; }

.HB1eCd-PLEiK-Tswv1b { background: rgb(246, 188, 93); color: rgb(34, 34, 34); }

.HB1eCd-PLEiK-Tswv1b-hSRGPd { color: rgb(6, 88, 181); }

.HB1eCd-PLEiK-GMvhG { background: rgb(204, 0, 0); color: rgb(255, 255, 255); }

.HB1eCd-PLEiK-GMvhG-hSRGPd { color: rgb(195, 217, 255); }

#docs-chrome-cover-container { width: 100%; z-index: 990; }

#docs-chrome-cover { height: 60px; }

#docs-transient-bar-container { left: 50%; position: absolute; top: 100%; width: 0px; }

.HB1eCd-JjiIAe-INgbqf-Ne3sFf { background-color: rgb(255, 255, 255); border-style: solid; border-color: rgb(153, 153, 153); border-image: initial; border-width: 0px 0px 1px; color: rgb(153, 153, 153); font-size: 28px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; position: absolute; text-align: center; }

.HB1eCd-r4nke-n0tgWb { margin-left: 17px; white-space: nowrap; }

.HB1eCd-r4nke-n0tgWb.HB1eCd-r4nke-TzA9Ye-Iqlsrf { margin-left: 12px; }

.HB1eCd-r4nke { display: inline-block; outline: none; }

.HB1eCd-r4nke-YPqjbf { border: 1px solid transparent; color: rgb(255, 255, 255); font-size: 18px; font-variant-ligatures: no-contextual; height: 20px; line-height: 22px; margin: 0px; min-width: 1px; padding: 2px 7px; visibility: hidden; border-radius: 2px !important; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-YPqjbf { font-size: 16px; }

.HB1eCd-r4nke-YPqjbf-V67aGc { font-size: 18px; font-variant-ligatures: no-contextual; line-height: 22px; margin: 0px; overflow: hidden; padding: 2px 8px; pointer-events: none; position: absolute; text-overflow: ellipsis; top: 0px; white-space: pre; z-index: 1; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-YPqjbf-V67aGc { font-size: 16px; }

.HB1eCd-r4nke-YPqjbf-V67aGc-SmKAyb { display: inline; line-height: 22px; }

.HB1eCd-r4nke-YPqjbf:hover { border-color: rgb(229, 229, 229); }

.HB1eCd-r4nke-YPqjbf:focus { appearance: none; box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; color: rgb(0, 0, 0); outline: none; border: 1px solid rgb(77, 144, 254) !important; }

.HB1eCd-r4nke-SmKAyb { color: rgb(51, 51, 51); font-size: 18px; max-width: 600px; margin: 2px 4px 1px 3px; overflow: hidden; text-overflow: ellipsis; white-space: pre; }

.HB1eCd-r4nke .HB1eCd-r4nke-NFS45c, .HB1eCd-r4nke-YPqjbf-V67aGc.HB1eCd-r4nke-NFS45c { color: rgb(119, 119, 119); font-style: italic; }

.HB1eCd-r4nke-m5SR9c { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 27px; width: auto; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-m5SR9c { padding-left: 6px; }

.HB1eCd-r4nke-m5SR9c-qnnXGd:hover .HB1eCd-r4nke { background-color: rgb(238, 238, 238); cursor: pointer; }

.HB1eCd-r4nke-m5SR9c .HB1eCd-a4fUwd-haAclf a { display: none; }

.HB1eCd-r4nke-m5SR9c:hover .HB1eCd-a4fUwd-haAclf a { display: inline-block; }

.HB1eCd-a4fUwd-haAclf { height: 21px; opacity: 0.6; padding-right: 9px; margin-top: 1px; vertical-align: top; width: 21px; }

.HB1eCd-a4fUwd-haAclf:hover { opacity: 0.9; }

.HB1eCd-NezmJd-KHwZ3c { vertical-align: top; }

.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-NezmJd-KHwZ3c > :not(.HB1eCd-ktSouf-uDEFge-haAclf) { display: none; }

.HB1eCd-NezmJd-Btuy5e-haAclf { padding: 0px 3px; vertical-align: top; }

.HB1eCd-NezmJd-Btuy5e .HB1eCd-Bz112c { display: block; height: 18px; margin: 3px; }

.HB1eCd-NezmJd-Btuy5e-haAclf .VIpgJd-bMcfAe, .HB1eCd-NezmJd-Btuy5e-haAclf .VIpgJd-Kb3HCc-LgbsSe { outline: none; }

.HB1eCd-NezmJd-Btuy5e { align-items: center; border-radius: 4px; color: rgb(95, 99, 104); cursor: pointer; display: flex; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; height: 24px; }

.HB1eCd-UMrnmb .HB1eCd-NezmJd-Btuy5e:hover, .HB1eCd-NezmJd-Btuy5e.VIpgJd-Kb3HCc-LgbsSe-XpnDCe, .HB1eCd-NezmJd-Btuy5e.VIpgJd-bMcfAe-XpnDCe, .VIpgJd-bMcfAe-XpnDCe .HB1eCd-NezmJd-Btuy5e { background-color: rgb(241, 243, 244); outline: none; }

.HB1eCd-UMrnmb .HB1eCd-NezmJd-Btuy5e:active, .HB1eCd-UMrnmb .HB1eCd-NezmJd-Btuy5e.HB1eCd-NezmJd-Btuy5e-gk6SMd { background-color: rgb(232, 240, 254); color: rgb(26, 115, 232); }

.HB1eCd-NezmJd-Btuy5e.VIpgJd-bMcfAe-OWB6Me { cursor: default; opacity: 0.38; background: none !important; }

.HB1eCd-NezmJd-Btuy5e.VIpgJd-bMcfAe-OWB6Me .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg") !important; }

.HB1eCd-NezmJd-KHwZ3c.HB1eCd-KHwZ3c-L6cTce-SfQLQb-QBLLGd { width: 0px; overflow: hidden; }

.HB1eCd-tlSJBe-hsovi-haAclf-n0tgWb { outline: none; vertical-align: top; }

.HB1eCd-Z0Arqf-uDEFge-haAclf { height: 29px; margin-top: 2px; vertical-align: top; padding-right: 2px; }

.S8Wip-QQhtn-TZk80d-IoWfhc-haAclf { display: inline-flex; }

.S8Wip-QQhtn-TZk80d-IoWfhc { background-color: rgb(26, 115, 232); border: 1px solid transparent; border-radius: 4px; box-sizing: border-box; color: rgb(255, 255, 255); cursor: default; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 13px; height: 21px; line-height: 21px; margin: 0px 8px 0px 0px; padding: 0px 5px 0px 4px; text-transform: uppercase; -webkit-font-smoothing: antialiased; }

.HB1eCd-Ujd07d-GQeX9e-VwQYGc-Btuy5e { margin: auto; }

.hXIJHe-S8Wip-QQhtn-TZk80d-IoWfhc { cursor: pointer; }

.HB1eCd-fTEazc-Btuy5e { border: 1px solid transparent; border-radius: 4px; box-sizing: border-box; cursor: pointer; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 12px; height: 20px; line-height: 15px; padding: 2px 8px; letter-spacing: 0.03em; }

.HB1eCd-NezmJd-Btuy5e-haAclf-L6cTce { padding: 0px; }

.HB1eCd-osrJF-Btuy5e-haAclf { vertical-align: middle; }

.HB1eCd-osrJF-Btuy5e { background-color: rgb(90, 90, 90); border-radius: 16px; color: white; font-size: 13px; padding: 0px 11px; height: 24px; line-height: 24px; }

#docs-dlp, #docs-activity-indicator { margin-left: 4px; outline: none; }

.HB1eCd-r4nke-ktSouf-V67aGc { outline: none; }

.HB1eCd-NezmJd-Btuy5e .HB1eCd-Bz112c-RJLb9c.HB1eCd-Bz112c-qknJed-AFZkUd { content: ""; }

.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-NezmJd-Btuy5e .HB1eCd-Bz112c-RJLb9c.HB1eCd-Bz112c-qknJed-AFZkUd { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

#docs-star.HB1eCd-NezmJd-Btuy5e:active { background-color: rgb(232, 234, 237); }

#docs-star.HB1eCd-NezmJd-Btuy5e:active .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); }

#docs-activity-indicator { padding-left: 4px; padding-top: 2px; }

#docs-dlp .HB1eCd-Bz112c-RJLb9c { opacity: 0.45; }

#docs-dlp:hover .HB1eCd-Bz112c-RJLb9c { opacity: 0.55; }

#docs-dlp, #docs-star, #docs-folder .HB1eCd-Bz112c { vertical-align: baseline; }

.HB1eCd-E90Ek-haAclf { margin-right: 6px; margin-top: 55px; vertical-align: top; font-size: 8px; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-E90Ek-haAclf { margin-top: calc(48px); }

.HB1eCd-NezmJd-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 0px 44px 0px 0px; position: absolute; right: 0px; text-align: right; top: 26px; vertical-align: middle; white-space: nowrap; box-sizing: border-box; }

.HB1eCd-E90Ek-haAclf.HB1eCd-E90Ek-Tswv1b { display: flex; position: absolute; right: 0px; top: 0px; }

.HB1eCd-NezmJd-LgbsSe { z-index: 1; }

#docs-docos-commentsbutton { margin-right: 9px; cursor: default; }

#docs-titlebar-save { text-align: center; }

#docs-docos-commentsbutton, #docs-titlebar-share-client-button div { height: 24px; padding-bottom: 3px; vertical-align: middle; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button div { height: 28px; margin-right: 8px; }

#docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button div.zAYgkb-Bz112c-LgbsSe { height: 32px; width: 32px; }

#docs-titlebar-share-client-button div.tk3N6e-LgbsSe { margin-right: 0px; }

.HB1eCd-NezmJd-c6xFrd .VIpgJd-xl07Ob-LgbsSe-j4gsHd { position: relative; top: 2px; vertical-align: baseline; }

.tk3N6e-O1htCb.VIpgJd-Kb3HCc-xl07Ob-LgbsSe > .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { text-align: left; }

.HB1eCd-loREFf { cursor: default; display: inline-block; font-size: 14px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 29px; margin-left: 52px; outline: none; position: relative; white-space: nowrap; }

.HB1eCd-loREFf .VIpgJd-bMcfAe { padding: 3px 7px 5px; margin-top: 2px; border: 1px solid transparent; outline: none; }

.HB1eCd-loREFf .VIpgJd-bMcfAe-ZmdkE { background: rgb(238, 238, 238); border-color: rgb(238, 238, 238); }

.HB1eCd-loREFf .VIpgJd-bMcfAe-FNFY6c { background: rgb(255, 255, 255); border-top: 1px solid rgba(0, 0, 0, 0.2); border-right: 1px solid rgba(0, 0, 0, 0.2); border-left: 1px solid rgba(0, 0, 0, 0.2); border-image: initial; border-bottom: none; box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; color: black; z-index: 1003; }

.HB1eCd-loREFf .VIpgJd-bMcfAe-OWB6Me { color: rgb(204, 204, 204); }

#docs-menubars { white-space: nowrap; }

#docs-editor-container { background: rgb(238, 238, 238); padding: 0px; }

#docs-editor { background: rgb(238, 238, 238); outline: none; }

#docs-editor.Kk7lMc-qnnXGd { width: calc(100% - 56px); }

.HB1eCd-w0UE8d-OWB6Me { color: rgb(153, 153, 153); cursor: text; }

.HB1eCd-ZYIfFd-V67aGc { display: none; }

.HB1eCd-r4nke-ktSouf-V67aGc { color: rgb(119, 119, 119); display: inline-block; margin-left: 14px; max-width: 250px; overflow: hidden; vertical-align: text-bottom; white-space: nowrap; }

.HB1eCd-r4nke-ktSouf-V67aGc-SfQLQb-Bz112c .HB1eCd-r4nke-ktSouf-V67aGc-fmcmS { max-width: calc(100% - 24px); }

.HB1eCd-r4nke-ktSouf-V67aGc-fmcmS { display: inline-block; max-width: 100%; overflow: hidden; text-overflow: ellipsis; vertical-align: text-bottom; white-space: nowrap; font-size: 14px; }

.HB1eCd-r4nke-ktSouf-V67aGc-fmcmS:hover, .HB1eCd-r4nke-ktSouf-V67aGc-fmcmS-XpnDCe { cursor: pointer; text-decoration: underline; }

.HB1eCd-r4nke-ktSouf-V67aGc-OWB6Me > .HB1eCd-r4nke-ktSouf-V67aGc-fmcmS:hover { cursor: auto; text-decoration: none; }

:not(.HB1eCd-r4nke-ktSouf-V67aGc-OWB6Me) > .HB1eCd-r4nke-ktSouf-V67aGc-fmcmS-hSRGPd { text-decoration: underline; }

.HB1eCd-HzV7m.HB1eCd-r4nke-ktSouf-V67aGc .HB1eCd-r4nke-ktSouf-V67aGc-Bz112c { cursor: pointer; margin: 0px 0px -1px 7px; opacity: 0.54; vertical-align: text-bottom; }

.HB1eCd-r4nke-ktSouf-V67aGc-fmcmS:empty + .HB1eCd-r4nke-ktSouf-V67aGc-Bz112c { display: none; }

.HB1eCd-r4nke-ktSouf-V67aGc-Ajmyi-wJBgYb { background-color: rgb(252, 228, 226); color: rgb(218, 54, 44); border-radius: 4px; margin-bottom: -5px; margin-left: 9px; padding: 5px; }

.HB1eCd-r4nke-ktSouf-V67aGc-Ajmyi-wJBgYb-LgbsSe { cursor: pointer; display: none; font-weight: bold; margin-left: 10px; outline: none; }

.HB1eCd-r4nke-ktSouf-V67aGc-Ajmyi-wJBgYb .HB1eCd-r4nke-ktSouf-V67aGc-Ajmyi-wJBgYb-LgbsSe { display: inline-block; }

.HB1eCd-r4nke-ktSouf-V67aGc-Ajmyi-wJBgYb-LgbsSe.VIpgJd-Kb3HCc-LgbsSe-OWB6Me { cursor: default; color: rgba(0, 0, 0, 0.26); }

#blob-notice-button { border: none; border-radius: 4px; background-color: rgb(252, 232, 230); color: rgb(197, 34, 31); cursor: pointer; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; margin: 0px 0px 0px 14px; outline: 0px; padding: 4px 8px; white-space: nowrap; }

.HB1eCd-Guievd-WqyaDf#blob-notice-button { border: 1px solid transparent; }

.S8Wip-QQhtn-zozyIf-u0pjoe-Ajmyi-wJBgYb-Bz112c, .S8Wip-QQhtn-GqqPG-u0pjoe-Ajmyi-wJBgYb-Bz112c { display: none; height: 14px; margin-left: -2px; margin-right: 2px; top: -1.5px; }

.HB1eCd-Iqlsrf-Sx9Kwc, .HB1eCd-DyVDA-ij8cu-Sx9Kwc { width: 340px; }

.HB1eCd-Iqlsrf-Sx9Kwc .XKSfm-Sx9Kwc-dI4VCc, .HB1eCd-DyVDA-ij8cu-Sx9Kwc .XKSfm-Sx9Kwc-dI4VCc { width: 300px; }

.HB1eCd-UMrnmb .HB1eCd-Iqlsrf-Sx9Kwc, .HB1eCd-UMrnmb .HB1eCd-DyVDA-ij8cu-Sx9Kwc { min-width: 312px; width: unset; }

.HB1eCd-UMrnmb .HB1eCd-Iqlsrf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { font-size: 12px; }

.HB1eCd-UMrnmb .HB1eCd-Iqlsrf-Sx9Kwc .XKSfm-Sx9Kwc-dI4VCc { width: 100%; }

#docs-help-anchor { left: 30%; position: absolute; }

#docs-help-anchor-right { right: 0px; position: absolute; }

.HB1eCd-AuE86-hSRGPd { color: rgb(34, 0, 204); cursor: pointer; text-decoration: underline; }

.HB1eCd-ynRLnc { position: absolute; left: -10000px; top: -10000px; }

.HB1eCd-ynRLnc-DmJKAe-cQYSPc { position: absolute; left: 0px; top: -1px; z-index: -2; opacity: 0; }

.VIpgJd-TUo6Hb-xJ5Hnf { z-index: 998; }

.VIpgJd-TUo6Hb { z-index: 1003; }

.VIpgJd-xl07Ob { z-index: 1003; }

#docs-menu-shield { background-color: rgb(255, 255, 255); position: absolute; z-index: 1004; }

.IyROMc-xl07Ob-ZYIfFd-bLicMb .VIpgJd-j7LFlb-PQTlnb-brjg8b { text-decoration: none; }

.IyROMc-xl07Ob-ZYIfFd-bLicMb .VIpgJd-j7LFlb-PQTlnb-hgDUwe { display: none; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-KEZkZ .HB1eCd-wckcKc { padding-left: 12px; color: rgb(154, 160, 166) !important; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-KEZkZ .IyROMc-j7LFlb { padding-right: 10px; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-GP8zAc .VIpgJd-j7LFlb.IyROMc-j7LFlb { padding-left: 16px; }

.VIpgJd-TzA9Ye-eEGnhe.HB1eCd-Bz112c.VIpgJd-j7LFlb-Bz112c { position: absolute; }

.VIpgJd-j7LFlb.IyROMc-j7LFlb { padding: 6px 10px 6px 30px; white-space: normal; }

.IyROMc-j7LFlb .VIpgJd-j7LFlb-V67aGc { padding-right: 6px; }

.IyROMc-j7LFlb .VIpgJd-j7LFlb-x29Bmf, .HB1eCd-UMrnmb .VIpgJd-j7LFlb .VIpgJd-j7LFlb-x29Bmf { float: right; padding: 0px 0px 0px 24px; position: relative; }

.VIpgJd-eKm5Fc .VIpgJd-j7LFlb-bN97Pc { margin-right: 42px; }

.HB1eCd-mZGCQb .VIpgJd-eKm5Fc-hFsbo, .IyROMc-j7LFlb .VIpgJd-eKm5Fc-hFsbo, .HB1eCd-UMrnmb .VIpgJd-j7LFlb .VIpgJd-eKm5Fc-hFsbo { margin-right: 4px; }

.XKSfm-Sx9Kwc-bN97Pc { font-size: 14px; }

#docs-hub-open-external-appbarbutton .R1gDOc-FNFY6c-HzdVzc-Bz112c-haAclf, #docs-hub-close-appbarbutton .R1gDOc-TvD9Pc-Bz112c-haAclf, .HB1eCd-Bz112c.VIpgJd-TzA9Ye-eEGnhe.R1gDOc-OMz1o-Bz112c-haAclf { height: 20px; outline: 0px; width: 20px; margin-top: 2px; }

.HB1eCd-MqDS2b-uoC0bf #docs-hub-open-external-appbarbutton .R1gDOc-FNFY6c-HzdVzc-Bz112c-haAclf, .HB1eCd-MqDS2b-uoC0bf #docs-hub-close-appbarbutton .R1gDOc-TvD9Pc-Bz112c-haAclf { height: 24px; left: 0px; top: 0px; width: 24px; }

#docs-hub-open-external-appbarbutton .R1gDOc-FNFY6c-HzdVzc-Bz112c-haAclf, #docs-hub-close-appbarbutton .R1gDOc-TvD9Pc-Bz112c-haAclf { position: relative; top: 1px; left: 1px; }

#docs-hub-open-external-appbarbutton, #docs-hub-close-appbarbutton { margin: 0px 0px 0px 2px; width: 32px; height: 32px; }

.HB1eCd-MqDS2b-uoC0bf #docs-hub-open-external-appbarbutton, .HB1eCd-MqDS2b-uoC0bf #docs-hub-close-appbarbutton { width: 36px; height: 36px; }

#docs-hub-open-external-appbarbutton:hover, #docs-hub-open-external-appbarbutton:focus, #docs-hub-close-appbarbutton:hover, #docs-hub-close-appbarbutton:focus { background-color: rgba(0, 0, 0, 0.06); }

input { font-family: inherit; }

.HB1eCd-RmniWd-Btuy5e { background-color: rgb(26, 115, 232); border-radius: 8px; color: rgb(255, 255, 255); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 500; height: 16px; letter-spacing: 0.3px; line-height: 16px; padding: 0px 6px; }

.HB1eCd-HzV7m #docs-branding-container { margin-top: 0px; width: 64px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c, .HB1eCd-HzV7m #docs-branding-container a, .HB1eCd-HzV7m #docs-branding-logo, .HB1eCd-HzV7m #docs-drive-logo { height: 40px; width: 40px; }

.HB1eCd-HzV7m #docs-branding-container a, .HB1eCd-HzV7m #docs-branding-container .HB1eCd-n7vHCb-l4eHX-di8rgd-hSRGPd { border-radius: 50%; margin: 4px 0px 4px 8px; padding: 8px; }

.HB1eCd-HzV7m #docs-branding-container a:focus { background-color: rgba(0, 0, 0, 0.06); outline: none; }

.HB1eCd-HzV7m #docs-menubar, .HB1eCd-HzV7m #docs-titlebar-container { margin-left: 64px; }

.HB1eCd-HzV7m .HB1eCd-r4nke-n0tgWb { margin-left: 0px; }

.HB1eCd-HzV7m #docs-folder:not(.HB1eCd-NezmJd-Btuy5e) { margin-top: 1px; }

.HB1eCd-HzV7m #docs-branding-container { background-color: inherit; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531.svg"); }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-TftRv { left: -20px; top: -4848px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-gvHUI { left: -20px; top: -320px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-TftRv-u2z5K { left: -22px; top: -9054px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-QymXn { left: -20px; top: -10248px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-QymXn-u2z5K { left: -26px; top: 0px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-zTETae, .HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-t02dhe, .HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-jdTLZc, .HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-ndfHFb { left: 0px; top: -11366px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-G1jlMc { left: 0px; top: -12142px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-G1jlMc-FMvwCe { left: 0px; top: -12938px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-G1jlMc-u2z5K { left: -20px; top: -11900px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-arrpzb { left: 0px; top: -5216px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-arrpzb-FMvwCe { left: 0px; top: -2180px; }

.HB1eCd-HzV7m .HB1eCd-n7vHCb-Bz112c-arrpzb-u2z5K { left: 0px; top: -6276px; }

.HB1eCd-HzV7m #docs-branding-container:not(.HB1eCd-n7vHCb-OQ09Xb-RCfa3e-OWB6Me):hover #docs-drive-logo { opacity: 0; }

.HB1eCd-HzV7m #docs-branding-container:not(.HB1eCd-n7vHCb-OQ09Xb-RCfa3e-OWB6Me):hover #docs-branding-logo { opacity: 1; }

.HB1eCd-HzV7m #docs-activity-indicator { padding-top: 3px; }

.HB1eCd-HzV7m .HB1eCd-NezmJd-KHwZ3c .tk3N6e-YhdZJc { vertical-align: top; }

.HB1eCd-HzV7m #docs-header #docs-titlebar { padding-top: 9px; }

.HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar { padding-top: calc(14px); }

.HB1eCd-HzV7m #docs-header #docs-titlebar-container { max-height: 33px; }

.HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-container { margin-left: 0px; max-height: none; }

.HB1eCd-HzV7m .HB1eCd-loREFf { height: 31px; }

.HB1eCd-HzV7m #docs-branding-container, .HB1eCd-HzV7m #docs-chrome-cover { height: 64px; }

.VIpgJd-INgbqf-LgbsSe, .VIpgJd-INgbqf-xl07Ob-LgbsSe { border-radius: 2px; user-select: none; background: 0px center; border-color: transparent; border-style: solid; border-width: 1px; outline: none; padding: 0px; height: 24px; color: rgb(68, 68, 68); line-height: 24px; list-style: none; text-decoration: none; vertical-align: middle; cursor: default; }

.VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border: 0px; vertical-align: top; }

.VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { margin: 0px; padding: 0px; }

.VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { padding: 0px 2px; }

.VIpgJd-INgbqf-LgbsSe-ZmdkE { padding: 0px; }

.VIpgJd-INgbqf-LgbsSe-auswjd, .VIpgJd-INgbqf-LgbsSe-barxie, .VIpgJd-INgbqf-LgbsSe-gk6SMd { color: rgb(34, 34, 34); padding: 0px; }

.VIpgJd-INgbqf-LgbsSe-ZmdkE, .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE { color: rgb(34, 34, 34); border-color: rgb(198, 198, 198) !important; }

.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { color: rgb(34, 34, 34); }

.VIpgJd-INgbqf-LgbsSe-ZmdkE, .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); }

.VIpgJd-INgbqf-LgbsSe-auswjd, .VIpgJd-INgbqf-xl07Ob-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(246, 246, 246); background-image: -webkit-linear-gradient(top, rgb(246, 246, 246), rgb(241, 241, 241)); border-color: rgb(198, 198, 198); }

.VIpgJd-INgbqf-LgbsSe-gk6SMd, .VIpgJd-INgbqf-LgbsSe-barxie, .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border-color: rgb(204, 204, 204); }

.VIpgJd-INgbqf-LgbsSe-OWB6Me, .VIpgJd-INgbqf-xl07Ob-LgbsSe-OWB6Me { opacity: 0.3; color: rgb(34, 34, 34) !important; }

.VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me, .VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { margin-right: 0px; }

.VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu, .VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { margin-left: 0px; }

.VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/ui/v1/disclosure/small-grey-disclosure-arrow-down.png") center center no-repeat; float: right; margin: 10px 2px 0px 3px; padding: 0px; opacity: 0.8; vertical-align: middle; width: 5px; height: 7px; }

.VIpgJd-INgbqf-hgDUwe { border-left: 1px solid rgb(204, 204, 204); height: 17px; line-height: normal; list-style: none; margin: 0px 2px; outline: none; overflow: hidden; padding: 0px; text-decoration: none; vertical-align: middle; width: 0px; }

.VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/ui/v1/disclosure/small-grey-disclosure-arrow-down.png") center center no-repeat; height: 11px; margin-top: 7px; width: 7px; transform: none; filter: none; }

.VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { padding: 0px; margin: 0px; }

.HB1eCd-HzV7m #docs-toolbar-wrapper { border-top: 1px solid rgb(224, 224, 224); border-bottom: 1px solid rgb(224, 224, 224); background: rgb(255, 255, 255); box-shadow: none; }

.HB1eCd-UMrnmb #docs-toolbar-wrapper { border-top: 1px solid rgb(218, 220, 224); border-bottom: 1px solid rgb(218, 220, 224); }

.HB1eCd-HzV7m #docs-side-toolbar { margin: 0px 21px 0px 0px; }

.HB1eCd-HzV7m.Kk7lMc-qnnXGd #docs-side-toolbar { margin: 0px 4px 0px 0px; }

.HB1eCd-HzV7m #docs-toolbar-wrapper, .HB1eCd-HzV7m #docs-equationtoolbar, .HB1eCd-HzV7m .HB1eCd-iqoopb-INgbqf { padding: 0px 21px 0px 22px; }

.HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-container { padding: 0px 21px 0px 24px; }

.HB1eCd-HzV7m #docs-equationtoolbar, .HB1eCd-HzV7m .HB1eCd-iqoopb-INgbqf { background: rgb(255, 255, 255); }

.HB1eCd-HzV7m #docs-equationtoolbar { border-top-width: 0px; border-bottom: 1px solid rgb(224, 224, 224); }

.HB1eCd-HzV7m.Kk7lMc-qnnXGd #docs-equationtoolbar { padding-right: 4px; }

.HB1eCd-UMrnmb #docs-equationtoolbar .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { padding-top: 0px; }

.HB1eCd-UMrnmb #docs-equationtoolbar .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { padding-top: 2px; }

#hide-equation-toolbar-button { float: right; }

#docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf { height: 26px; line-height: 26px; }

#docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf::placeholder { line-height: 26px; }

#docs-omnibox-toolbar .HB1eCd-QbdDtf-h0T7hb { margin: 6px 4px 6px 1px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf, .HB1eCd-UMrnmb #docs-toolbar { min-height: 38px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe, .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe { box-shadow: none; background-color: rgb(255, 255, 255); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-WTFKld-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m.xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-ZmdkE { box-shadow: none; background-color: rgba(0, 0, 0, 0.06); background-image: none; border-radius: 2px; border-width: 1px; cursor: pointer; border-color: transparent !important; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-WTFKld-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-PimBUc-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-LgbsSe-hgDUwe-sM5MNb, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE .HB1eCd-UMrnmb .HB1eCd-HzV7m.xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-ZmdkE { background-color: rgb(241, 243, 244); }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-auswjd, .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie, .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-gk6SMd, .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-LgbsSe-auswjd, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-auswjd, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { box-shadow: none; background-color: rgba(0, 0, 0, 0.12); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m.xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd { box-shadow: none; background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-gk6SMd, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m.xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd { background-color: rgb(232, 240, 254); color: rgb(26, 115, 232); }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe { margin: 3px 1px 0px; height: 26px; line-height: 26px; color: rgba(0, 0, 0, 0.7); }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { height: 26px; min-width: 26px; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { min-width: 26px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie + .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie { border-left: 1px solid rgb(204, 204, 204); border-top-left-radius: 2px; border-bottom-left-radius: 2px; margin-left: 1px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie + .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .HB1eCd-HzV7m .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie + .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie.VIpgJd-INgbqf-LgbsSe-ZmdkE .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { margin-left: 0px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe .HB1eCd-Bz112c { opacity: 0.54; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { opacity: 1; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-ZmdkE .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-gk6SMd .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-auswjd .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-gk6SMd .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-barxie .HB1eCd-Bz112c, .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c .HB1eCd-Bz112c { opacity: 0.87; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-ZmdkE .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-gk6SMd .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-auswjd .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-gk6SMd .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-barxie .HB1eCd-Bz112c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c .HB1eCd-Bz112c { opacity: 1; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .HB1eCd-UMrnmb .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { height: 24px; min-width: 24px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-LgbsSe .HB1eCd-Bz112c { margin: 0px 0px 1px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-LgbsSe.HB1eCd-Bz112c-INgbqf-LgbsSe-SfQLQb-fmcmS .HB1eCd-Bz112c-INgbqf-LgbsSe-SfQLQb-fmcmS-Bz112c-haAclf { margin-right: 4px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-xl07Ob-LgbsSe.HB1eCd-vJX8Jf .HB1eCd-Bz112c { margin-top: 1px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-hgDUwe.VIpgJd-TzA9Ye-eEGnhe { border-left: 1px solid rgb(224, 224, 224); margin: 0px 3px; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-purZT-hgDUwe + div.VIpgJd-INgbqf-LgbsSe, .HB1eCd-HzV7m .HB1eCd-INgbqf-purZT-hgDUwe + div.VIpgJd-INgbqf-xl07Ob-LgbsSe { margin-left: 1px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-hgDUwe.VIpgJd-TzA9Ye-eEGnhe { border-left: 1px solid rgb(218, 220, 224); margin: 9px 4px; height: 20px; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu.VIpgJd-TzA9Ye-eEGnhe { margin-right: 0px; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-TzA9Ye-eEGnhe { margin-left: 0px; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.HB1eCd-INgbqf-LgbsSe-DIdRlc-WTFKld-ZmdkE, .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu + .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe + .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me { border-left-color: rgba(0, 0, 0, 0.12) !important; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.HB1eCd-INgbqf-LgbsSe-DIdRlc-WTFKld-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu + .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe + .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me { border-left-color: rgb(241, 243, 244) !important; }

.HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe { margin-right: 3px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-HzV7m .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-HzV7m .VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd { margin-top: 10px; }

.HB1eCd-UMrnmb .HB1eCd-UMrnmb-hFsbo .HB1eCd-Bz112c { margin: 0px; }

.HB1eCd-HzV7m .VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { margin-top: 8px; }

.HB1eCd-UMrnmb .HB1eCd-UMrnmb-hFsbo.VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .HB1eCd-INgbqf-DIdRlc-t0O6ic-LgbsSe .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .HB1eCd-UMrnmb-hFsbo.VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd { background: none; margin: 0px -1px 0px -3px; width: 13px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { margin-right: -1px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-LgbsSe, .HB1eCd-UMrnmb .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .VIpgJd-INgbqf-yiAvpe-LgbsSe, .HB1eCd-UMrnmb #docs-equationtoolbar .VIpgJd-INgbqf-LgbsSe, .HB1eCd-UMrnmb #docs-equationtoolbar .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf { height: 24px; line-height: 24px; margin: 6px 1px; top: 0px; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .VIpgJd-INgbqf-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-OWB6Me { cursor: inherit; opacity: 0.38; color: rgb(95, 99, 104) !important; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { color: rgba(0, 0, 0, 0.7); box-sizing: border-box; height: 20px !important; width: 48px !important; }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf::selection { background-color: rgb(232, 240, 254); }

.HB1eCd-UMrnmb .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf:focus { border-radius: 4px; padding: 0px 7px; border: 2px solid rgb(26, 115, 232) !important; }

.HB1eCd-HzV7m .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge { height: 20px; border-bottom-color: transparent; forced-color-adjust: none; }

.HB1eCd-HzV7m .HB1eCd-vJX8Jf .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge { bottom: 0px; }

.HB1eCd-HzV7m.HB1eCd-INgbqf-z5C9Gb-VCkuzd { border: 0px; box-shadow: rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 3px 1px -2px, rgba(0, 0, 0, 0.2) 0px 1px 5px 0px; border-radius: 2px; }

.HB1eCd-HzV7m.HB1eCd-INgbqf-z5C9Gb-VCkuzd .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG, .HB1eCd-HzV7m.HB1eCd-INgbqf-z5C9Gb-VCkuzd .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { border-color: transparent; }

.HB1eCd-HzV7m.HB1eCd-INgbqf-z5C9Gb-INgbqf { background: rgb(255, 255, 255); border-radius: 2px; padding: 0px 4px; }

.HB1eCd-UMrnmb .HB1eCd-INgbqf-z5C9Gb-VCkuzd { border-radius: 4px; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb .HB1eCd-INgbqf-z5C9Gb-INgbqf { border-radius: 4px; }

::-webkit-scrollbar { height: 16px; overflow: visible; width: 16px; }

::-webkit-scrollbar-button { height: 0px; width: 0px; }

::-webkit-scrollbar-track { background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 0px 0px 0px 4px; }

::-webkit-scrollbar-track:horizontal { border-width: 4px 0px 0px; }

::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.1) 1px 0px 0px inset; }

::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 0px inset; }

::-webkit-scrollbar-track:active { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.2) 1px 0px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(255, 255, 255, 0.2) 0px 1px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:active { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.25) 1px 0px 0px inset, rgba(255, 255, 255, 0.15) -1px 0px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(255, 255, 255, 0.25) 0px 1px 0px inset, rgba(255, 255, 255, 0.15) 0px -1px 0px inset; }

::-webkit-scrollbar-thumb { background-color: rgba(0, 0, 0, 0.2); background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 1px 1px 1px 6px; min-height: 28px; padding: 100px 0px 0px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

::-webkit-scrollbar-thumb:horizontal { border-width: 6px 1px 1px; padding: 0px 0px 0px 100px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

::-webkit-scrollbar-thumb:hover { background-color: rgba(0, 0, 0, 0.4); box-shadow: rgba(0, 0, 0, 0.25) 1px 1px 1px inset; }

::-webkit-scrollbar-thumb:active { background-color: rgba(0, 0, 0, 0.5); box-shadow: rgba(0, 0, 0, 0.35) 1px 1px 3px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb { background-color: rgba(255, 255, 255, 0.3); box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) 0px -1px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:horizontal { box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) -1px 0px 0px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:hover { background-color: rgba(255, 255, 255, 0.6); box-shadow: rgba(255, 255, 255, 0.37) 1px 1px 1px inset; }

.tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:active { background-color: rgba(255, 255, 255, 0.75); box-shadow: rgba(255, 255, 255, 0.5) 1px 1px 3px inset; }

.tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track { border-width: 0px 1px 0px 6px; }

.tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track:horizontal { border-width: 6px 0px 1px; }

.tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.035); box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px -1px 0px inset; }

.tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.07); box-shadow: rgba(255, 255, 255, 0.25) 1px 1px 0px inset, rgba(255, 255, 255, 0.15) -1px -1px 0px inset; }

.tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-thumb { border-width: 0px 1px 0px 6px; }

.tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-thumb:horizontal { border-width: 6px 0px 1px; }

::-webkit-scrollbar-corner { background: transparent; }

body::-webkit-scrollbar-track-piece { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 0px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

body::-webkit-scrollbar-track-piece:horizontal { border-width: 3px 0px 0px; box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

body::-webkit-scrollbar-thumb { border-width: 1px 1px 1px 5px; }

body::-webkit-scrollbar-thumb:horizontal { border-width: 5px 1px 1px; }

body::-webkit-scrollbar-corner { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 3px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset; }

.tk3N6e-LgbsSe { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.VIpgJd-INgbqf-LgbsSe, .VIpgJd-INgbqf-xl07Ob-LgbsSe { font-weight: 500; font-size: 12px; }

.HB1eCd-UMrnmb #docs-editor, .HB1eCd-UMrnmb #docs-editor-container { background: rgb(248, 249, 250); }

.HB1eCd-MqDS2b-uoC0bf #docs-editor, .HB1eCd-MqDS2b-uoC0bf #docs-editor-container { background: rgb(249, 251, 253); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-R1gDOc #docs-editor-container { background: rgb(255, 255, 255); }

.VIpgJd-AznF2e { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { font-weight: 400; }

.XKSfm-Sx9Kwc-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.tk3N6e-F79BRe .VIpgJd-VgwJlc-PBWx0c, .tk3N6e-eLJrl { font-weight: 500; }

.tk3N6e-rugWtd-xGWjg, .tk3N6e-rugWtd-xGWjg:hover { font-weight: 500; }

.tk3N6e-suEOdc { font-weight: 500; font-size: 12px; }

.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc, .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { border-color: rgb(218, 220, 224) transparent; }

@media (forced-colors: active) {
  .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd.HB1eCd-EfADOe-VCkuzd { border: 1px solid canvastext; }
  .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG, .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc, .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border-color: canvastext canvas; }
  @supports (forced-color-adjust: none) {
  .tk3N6e-suEOdc-jQ8oHc, .tk3N6e-suEOdc-ez0xG, .HB1eCd-UMrnmb-EfADOe .tk3N6e-VCkuzd-jQ8oHc, .HB1eCd-UMrnmb-EfADOe .tk3N6e-VCkuzd-ez0xG { forced-color-adjust: none; }
  .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc { border-color: canvastext transparent; }
  .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { border-color: canvas transparent; }
  .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd.tk3N6e-VCkuzd-EfADOe.HB1eCd-EfADOe-VCkuzd .tk3N6e-VCkuzd-hFsbo-hUbt4d.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border-color: canvastext transparent; }
}
}

.IyROMc-t6O8cf-r4nke-haAclf, .IyROMc-w3KqTd-r4nke-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb .HB1eCd-E90Ek-haAclf { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb .HB1eCd-tCYPLb-LkdAo, .HB1eCd-UMrnmb .HB1eCd-tCYPLb-DbqQVb, .HB1eCd-UMrnmb .HB1eCd-jEqmyf-oPu43, .HB1eCd-UMrnmb .pD2Zae-k6D2ve-cXXICe-LYNcwc { background-color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb .HB1eCd-tCYPLb-i5vt6e, .HB1eCd-UMrnmb .HB1eCd-jEqmyf-VtOx3e, .HB1eCd-UMrnmb .HB1eCd-bwj4ec-VtOx3e { border-color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb .HB1eCd-tCYPLb-DbqQVb { height: 24px; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); cursor: pointer; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-QDgCrf { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; cursor: default; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); cursor: pointer; border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-QDgCrf, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-QDgCrf, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-QDgCrf { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; cursor: default; border: 1px solid rgb(241, 243, 244) !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:hover, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:focus, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:focus, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { border: 1px solid highlight; }
}

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:hover:focus, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:active, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc button:focus:active, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc button[disabled], .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; border: 1px solid rgb(241, 243, 244) !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); border: 1px solid transparent !important; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:hover, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:focus, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:hover:focus, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:active, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:focus:active, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc[disabled], .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-LgbsSe, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc button, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc { cursor: pointer; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-LgbsSe.VIpgJd-Kb3HCc-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc button[disabled], .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc[disabled], .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { cursor: default; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .tk3N6e-y4JFTd, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-y4JFTd, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(60, 64, 67); padding: 1px 8px; font-size: 14px; height: 36px; margin: 8px 0px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc textarea.tk3N6e-y4JFTd { min-height: 36px; height: unset; padding: 7px 8px; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc textarea.tk3N6e-y4JFTd { min-height: 52px; max-height: 52px; min-width: 100%; height: unset; padding: 7px 8px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb .HB1eCd-HzV7m-VCkuzd .tk3N6e-y4JFTd:focus { border: 2px solid rgb(26, 115, 232); box-shadow: none; padding: 0px 7px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc textarea.tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc textarea.tk3N6e-y4JFTd:focus { padding: 6px 7px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { background-color: transparent; border-radius: 50%; cursor: pointer; line-height: 18px; text-align: center; color: rgb(95, 99, 104); }

.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: rgb(232, 234, 237); outline: none; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { color: canvastext; }
  .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: highlight; color: highlighttext; }
}

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd.EX2EHc-cwdWJf-rygyx { margin: 0px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc.jcJzye-dZ8yzd-fFW7wc, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF.tk3N6e-VCkuzd, .HB1eCd-UMrnmb .HB1eCd-Yygnk-uDEFge-V68bde.tk3N6e-VCkuzd { background: rgb(255, 255, 255); border: 1px solid transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; position: absolute; z-index: 1003; padding: 24px; }

.HB1eCd-UMrnmb .fFW7wc.XKSfm-Sx9Kwc { padding: 0px; z-index: 1201; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc.jcJzye-dZ8yzd-fFW7wc, .HB1eCd-UMrnmb .XKSfm-Sx9Kwc-bN97Pc, .HB1eCd-UMrnmb #docs-offline-optinpromo-description, .HB1eCd-UMrnmb #docs-offline-optinpromo-learn-more-container { color: rgb(60, 64, 67); }

.HB1eCd-UMrnmb #docs-offline-optinpromo-title { border-bottom: none; padding: 24px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc-r4nke-fmcmS, .HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-r4nke-fmcmS { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 22px; font-weight: 400; line-height: 28px; }

.HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd { display: flex; flex-direction: row-reverse; }

.HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-McfNlf-c6xFrd { margin-top: 24px; }

.HB1eCd-UMrnmb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe { cursor: pointer; margin-left: 16px; margin-right: 0px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc-c6xFrd, .HB1eCd-UMrnmb .HB1eCd-NRdnKf-c6xFrd { display: flex; justify-content: flex-end; margin-top: 24px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc-c6xFrd button { margin: 0px 0px 0px 12px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc-c6xFrd button:first-child { margin-left: 0px; }

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { position: relative; }

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-fmcmS { display: inline-block; max-width: calc(100% - 32px); min-width: 200px; }

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc { background-color: transparent; border-radius: 50%; cursor: pointer; height: 18px; line-height: 18px; padding: 7px; right: 0px; text-align: center; top: -3px; width: 18px; }

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:hover { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: rgb(232, 234, 237); outline: none; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:focus { border: 1px solid highlight; padding: 6px; }
}

.HB1eCd-UMrnmb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc::after { position: relative; right: 0px; top: 0px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { height: 22px; width: 22px; border-radius: 50%; border: 1px solid rgb(218, 220, 224); margin: 0px; outline: none; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { padding: 6px 0px 6px 6px; }

.HB1eCd-UMrnmb div.VIpgJd-TUo6Hb-xJ5Hnf, .HB1eCd-UMrnmb div.XKSfm-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); left: 0px; position: absolute; top: 0px; z-index: 998; opacity: 0.6 !important; }

.HB1eCd-UMrnmb ::-webkit-scrollbar-track { box-shadow: none; margin: 0px 4px; }

.HB1eCd-UMrnmb ::-webkit-scrollbar-track:hover { box-shadow: none; background: none; }

.HB1eCd-UMrnmb ::-webkit-scrollbar-thumb { border-style: solid; border-color: transparent; border-width: 4px; background-color: rgb(218, 220, 224); border-radius: 8px; box-shadow: none; }

.HB1eCd-UMrnmb ::-webkit-scrollbar-thumb:hover { background-color: rgb(128, 134, 139); }

.HB1eCd-UMrnmb ::-webkit-scrollbar-thumb:active { background-color: rgb(95, 99, 104); }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; cursor: pointer; padding: 8px 6px 8px 8px; align-items: center; background: none; color: rgb(60, 64, 67); display: inline-flex; justify-content: space-between; outline: none; position: relative; width: unset; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { color: rgb(95, 99, 104); opacity: 0.38; cursor: default; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active { background-color: rgb(255, 255, 255); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { background-color: rgba(60, 64, 67, 0.04); border: 1px solid rgb(218, 220, 224); box-shadow: none; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { background-color: rgba(60, 64, 67, 0.06); border: 1px solid rgb(218, 220, 224); }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { border: 1px solid highlight; }
}

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.04); border: 1px solid transparent; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.06); }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.08); }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { border: 1px solid rgb(218, 220, 224); box-shadow: none; cursor: default; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { box-sizing: border-box; color: rgb(32, 33, 36); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; height: 20px; line-height: 20px; max-width: 100%; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { color: rgb(95, 99, 104); opacity: 0.38; cursor: default; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg") -48px -12142px no-repeat; height: 18px; width: 18px; border: none; margin-top: 0px; position: relative; right: 0px; top: 0px; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { opacity: 0.38; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active { border: 1px solid rgb(218, 220, 224); cursor: default; box-shadow: none; }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { transform: rotate(180deg); }

.HB1eCd-UMrnmb .XKSfm-Sx9Kwc .tk3N6e-Ru3Ixf-OWB6Me .tk3N6e-Ru3Ixf-V67aGc { color: rgb(95, 99, 104); opacity: 0.38; cursor: default; }

.HB1eCd-UMrnmb .euCgFf-X3SwIb-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; }

.HB1eCd-UMrnmb .euCgFf-CJXtmf-Sx9Kwc .euCgFf-X3SwIb-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb .euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd { height: 40px; padding: 0px 16px; }

.HB1eCd-UMrnmb .euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd > span { display: flex; padding-top: 4px; }

.HB1eCd-UMrnmb .euCgFf-PLEiK-Bz112c { margin-right: 8px; }

.HB1eCd-UMrnmb .euCgFf-PLEiK-hSRGPd, .HB1eCd-UMrnmb .euCgFf-PLEiK-hSRGPd:visited { color: rgb(26, 115, 232); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 16px; margin-left: 80px; }

.HB1eCd-UMrnmb .euCgFf-PLEiK-hSRGPd:hover, .HB1eCd-UMrnmb .euCgFf-PLEiK-hSRGPd:active { color: rgb(24, 90, 188); }

.HB1eCd-UMrnmb .euCgFf-PLEiK-hSRGPd:disabled { color: rgb(26, 115, 232); }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; background: rgb(194, 231, 255); color: rgb(0, 29, 53); }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe-OWB6Me, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; background: rgb(228, 228, 228); color: rgb(31, 31, 31); cursor: default; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe:focus, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:focus { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; color: rgb(0, 29, 53); background: rgb(171, 207, 231); box-shadow: none; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; color: rgb(0, 29, 53); background: rgb(178, 215, 239); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 1px 3px 1px; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE:focus, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE:focus { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; color: rgb(0, 29, 53); background: rgb(171, 207, 231); box-shadow: none; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-auswjd, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-barxie, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; color: rgb(0, 29, 53); background: rgb(150, 186, 210); }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .tk3N6e-LgbsSe .zAYgkb-LgbsSe-Bz112c { margin: 0px 8px 1px -8px; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe:focus, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE:focus, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-auswjd, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-barxie { border-bottom-right-radius: 0px; border-top-right-radius: 0px; padding: 10px 8px 10px 24px; margin-right: 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-DIdRlc-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE:focus, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE:focus { box-shadow: none; }

.HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:focus, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE:focus, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd { border-bottom-left-radius: 0px; border-left: 1px solid rgb(255, 255, 255); border-top-left-radius: 0px; padding-left: 0px; padding-right: 8px; margin-left: -1px; margin-right: 8px; min-width: 34px; width: 34px; }

.HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { opacity: 0.62; }

.HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd.VIpgJd-TzA9Ye-eEGnhe, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd.VIpgJd-TzA9Ye-eEGnhe { top: 18px; right: 12px; }

#docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe, #docs-titlebar-share-client-button .tk3N6e-LgbsSe-OWB6Me.zAYgkb-Bz112c-LgbsSe, #docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe.tk3N6e-LgbsSe-ZmdkE, #docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe.tk3N6e-LgbsSe-ZmdkE:focus, #docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe.tk3N6e-LgbsSe-auswjd, #docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe.tk3N6e-LgbsSe-XpnDCe { border-radius: 100%; padding: 10px; }

#docs-titlebar-share-client-button .tk3N6e-LgbsSe.zAYgkb-Bz112c-LgbsSe .zAYgkb-LgbsSe-Bz112c { margin: 0px 0px 2px; padding-right: 1px; }

.HB1eCd-MqDS2b-uoC0bf #docs-titlebar-share-client-button .zAYgkb-ti6hGc-b3rLgd::after, .HB1eCd-MqDS2b-uoC0bf #scb-quick-actions-menu-button .zAYgkb-ti6hGc-b3rLgd::after { background-color: rgb(11, 87, 208); border-radius: calc(5px); content: ""; min-height: 10px; min-width: 10px; outline: rgb(249, 251, 253) solid 2px; position: absolute; right: 0px; top: 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-header:not(.HB1eCd-R1gDOc-UU3Zxb) .HB1eCd-NezmJd-c6xFrd { background: rgb(249, 251, 253); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-docos-commentsbutton { margin-right: 6px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-docos-commentsbutton .HB1eCd-wvGCSb-Pqjfme-Btuy5e { background: rgb(11, 87, 208); font-family: "Google Sans", Roboto, sans-serif; letter-spacing: 0.25px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke-YPqjbf { background: none; padding: 1px 6px; color: rgb(249, 251, 253); border-radius: 4px !important; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-R1gDOc .HB1eCd-r4nke-YPqjbf { padding-top: 2px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke-YPqjbf-V67aGc { padding-left: 7px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-YPqjbf { color: rgb(255, 255, 255); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke .HB1eCd-r4nke-NFS45c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke-YPqjbf-V67aGc.HB1eCd-r4nke-NFS45c { color: rgb(68, 71, 70); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke-YPqjbf:focus { color: rgb(31, 31, 31); margin: 0px -1px; border-color: rgb(11, 87, 208) !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-r4nke-YPqjbf:hover { border-color: rgb(116, 119, 117); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e:active { color: rgb(95, 99, 104); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e.HB1eCd-NezmJd-Btuy5e-gk6SMd { background-color: rgb(225, 227, 230); color: rgb(95, 99, 104); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e .HB1eCd-ktSouf-uDEFge-Bz112c { border-radius: 50%; font-family: "Google Sans", Roboto, sans-serif; height: 28px; justify-content: center; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e:hover, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e .HB1eCd-ktSouf-uDEFge-Bz112c:hover { background-color: rgb(232, 235, 238); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e:active, .HB1eCd-MqDS2b-uoC0bf #docs-star.HB1eCd-NezmJd-Btuy5e:active, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e:focus, .HB1eCd-MqDS2b-uoC0bf .VIpgJd-bMcfAe-XpnDCe .HB1eCd-NezmJd-Btuy5e .HB1eCd-ktSouf-uDEFge-Bz112c, .HB1eCd-MqDS2b-uoC0bf .VIpgJd-bMcfAe-auswjd .HB1eCd-NezmJd-Btuy5e .HB1eCd-ktSouf-uDEFge-Bz112c { background-color: rgb(225, 227, 230); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e.HB1eCd-ktSouf-uDEFge:hover, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e.HB1eCd-ktSouf-uDEFge:active, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e.HB1eCd-ktSouf-uDEFge:focus, .HB1eCd-MqDS2b-uoC0bf .VIpgJd-bMcfAe-XpnDCe .HB1eCd-NezmJd-Btuy5e.HB1eCd-ktSouf-uDEFge, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e-gk6SMd.HB1eCd-ktSouf-uDEFge { background-color: transparent; }

.HB1eCd-MqDS2b-uoC0bf #docs-star.HB1eCd-NezmJd-Btuy5e:active .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e-haAclf { padding: 0px 2px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-Btuy5e .HB1eCd-Bz112c { height: 20px; width: 20px; margin: 4px; }

.HB1eCd-MqDS2b-uoC0bf #docs-star .HB1eCd-Bz112c-RJLb9c { margin-top: -1px; }

.HB1eCd-MqDS2b-uoC0bf #docs-header { height: 32px !important; }

.HB1eCd-MqDS2b-uoC0bf #docs-header.HB1eCd-R1gDOc-UU3Zxb { height: 55px !important; }

.HB1eCd-NezmJd-qAWA2#docs-header { height: 59px !important; }

#docs-header .HB1eCd-NezmJd-qAWA2#docs-titlebar-container { align-items: center; display: flex; height: 59px; max-height: 59px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-NezmJd-qAWA2#docs-titlebar-container #docs-titlebar { height: auto; padding-top: 12px; }

.HB1eCd-MqDS2b-uoC0bf #docs-menubars { margin-top: -6px; transition-duration: 100ms; height: auto !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header .HB1eCd-NezmJd-c6xFrd { height: 60px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header .HB1eCd-NezmJd-c6xFrd.HB1eCd-NezmJd-c6xFrd-nUpftc-WAutxc { height: 58px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-NezmJd-c6xFrd-nUpftc-WAutxc .HB1eCd-E90Ek-haAclf { margin-top: 50px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header #docs-titlebar { padding-top: 8px; }

.HB1eCd-MqDS2b-uoC0bf #docs-chrome.HB1eCd-R1gDOc-NMrWyd { border-color: transparent; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m .HB1eCd-R1gDOc-UU3Zxb#docs-header #docs-titlebar { height: 100%; padding-top: 0px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-n0tgWb { align-items: center; display: flex; height: 100%; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-NezmJd-c6xFrd { height: 100%; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button .tk3N6e-LgbsSe:not(.zAYgkb-Bz112c-LgbsSe) { padding: 8px 24px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button .tk3N6e-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-ZmdkE:focus, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button .tk3N6e-LgbsSe.tk3N6e-LgbsSe-auswjd { height: 36px; }

.HB1eCd-MqDS2b-uoC0bf #docs-header.HB1eCd-R1gDOc-UU3Zxb #docs-titlebar-share-client-button div.zAYgkb-Bz112c-LgbsSe { height: 36px; width: 36px; }

.HB1eCd-MqDS2b-uoC0bf #docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-YPqjbf { padding-top: 2px; font-size: 18px; }

.HB1eCd-MqDS2b-uoC0bf #docs-header.HB1eCd-R1gDOc-UU3Zxb .HB1eCd-r4nke-YPqjbf-V67aGc { font-size: 18px; top: 1px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-HzV7m #docs-toolbar-wrapper { background-color: rgb(237, 242, 250); border: none; border-radius: 24px; font-family: "Google Sans", Roboto, sans-serif; margin: 6px 16px 8px; min-height: 40px; padding: 0px 8px; -webkit-font-smoothing: antialiased; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-INgbqf-z5C9Gb-INgbqf, .HB1eCd-MqDS2b-uoC0bf .xih9X-nEeMgc { background-color: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { height: 28px; min-width: 28px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf.HB1eCd-UMrnmb #docs-toolbar-wrapper, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf #docs-align-palette, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf #docs-align-palette .VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .HB1eCd-INgbqf-z5C9Gb-INgbqf { background: rgb(243, 246, 252); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-O1htCb, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe { border-radius: 4px; height: 28px; line-height: 28px; margin: 5px 1px; min-width: 28px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe { border-radius: 4px; line-height: 28px; margin: 5px 1px; min-width: 28px; }

.HB1eCd-MqDS2b-uoC0bf #docs-equationtoolbar .VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #docs-equationtoolbar .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf { border-radius: 4px; height: 28px; line-height: 28px; margin: 5px 1px; min-width: 28px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .xih9X-nEeMgc .VIpgJd-INgbqf-xl07Ob-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #docs-align-palette .VIpgJd-INgbqf-LgbsSe { background-color: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .lUepf-nEeMgc .VIpgJd-nEeMgc-eEDwDf-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-INgbqf-nJjxad-Dd6Aae.VIpgJd-INgbqf-yiAvpe-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf .xih9X-nEeMgc .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb #docs-align-palette .VIpgJd-INgbqf-LgbsSe-ZmdkE { background-color: rgba(68, 71, 70, 0.08); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe { height: 26px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe:focus, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe-auswjd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-auswjd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe:focus, .HB1eCd-MqDS2b-uoC0bf .xih9X-nEeMgc .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(68, 71, 70, 0.12); color: rgb(68, 71, 70); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .lUepf-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb #docs-align-palette .VIpgJd-INgbqf-LgbsSe-barxie { background-color: rgb(211, 227, 253); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .lUepf-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf #docs-align-palette .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .lUepf-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .xih9X-nEeMgc .VIpgJd-nEeMgc-eEDwDf-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye #docs-align-palette .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(12%) sepia(17%) saturate(6039%) hue-rotate(199deg) brightness(93%) contrast(106%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae.VIpgJd-INgbqf-yiAvpe-LgbsSe { border-radius: 4px; border: 1px solid rgb(116, 119, 117) !important; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae.VIpgJd-INgbqf-yiAvpe-LgbsSe-ZmdkE { border: 1px solid rgb(31, 31, 31) !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c { border-radius: 4px; margin: 0px; border: 2px solid rgb(11, 87, 208) !important; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae.VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c { border-radius: 4px; border: 2px solid rgb(11, 87, 208) !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { color: rgb(68, 71, 70); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf:focus { box-shadow: none; padding: 0px 4px; background: transparent; border: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { color: rgb(68, 71, 70); padding: 1px 4px; font-family: "Google Sans", Roboto, sans-serif !important; font-size: 14px !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf:focus, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { color: rgb(31, 31, 31); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-ZmdkE .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { border-right: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-SmKAyb-Q4BLdf { margin: 0px 4px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-UMrnmb-hFsbo.VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd { margin-right: 2px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { margin-right: 4px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd .HB1eCd-Bz112c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd .HB1eCd-Bz112c { height: 18px; width: 18px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c .VIpgJd-INgbqf-yiAvpe-LgbsSe-j4gsHd .HB1eCd-Bz112c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-O1htCb.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd .HB1eCd-Bz112c { margin-bottom: 3px; transform: rotateX(180deg); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-HzV7m .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me { margin-left: 0px; border-color: transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-LgbsSe-DIdRlc-LK5yu { margin-right: 0px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-LgbsSe-DIdRlc-qwU8Me.VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { background-color: rgb(211, 227, 253); }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae { width: 32px !important; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { margin: -1px -1px -1px 0px; width: 32px !important; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeIncrement.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-JIbuQc-LgbsSe.VIpgJd-INgbqf-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #fontSizeDecrement.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-JIbuQc-LgbsSe.VIpgJd-INgbqf-LgbsSe { border: none; border-radius: 4px; height: 24px; width: 24px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-JIbuQc-LgbsSe .HB1eCd-Bz112c { margin: 2px 0px 0px 1px; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae { margin: 0px 3px; border-color: transparent !important; }

.HB1eCd-MqDS2b-uoC0bf #fontSizeSelect.HB1eCd-sLO9V-SxQuSe-WXLSre-TLR7cb-Dd6Aae.VIpgJd-INgbqf-yiAvpe-LgbsSe-FNFY6c { margin: 0px 2px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-h0T7hb { margin: 3px 2px 6px 1px; padding: 2px 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf { background: white; border-radius: 28px; color: rgb(31, 31, 31); height: 28px; line-height: 32px; padding-left: 16px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd[aria-expanded="true"] { border-bottom: rgb(225, 227, 225); border-radius: 8px 8px 0px 0px; padding-left: 16px; }

.HB1eCd-MqDS2b-uoC0bf #docs-toolbar.VIpgJd-INgbqf { padding-left: 2px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-Bz112c { margin: 5px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-oKdM2c-Bz112c { margin-top: 1px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf::placeholder { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf::selection { background-color: rgb(211, 227, 253); }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-fmcmS-LgbsSe .VIpgJd-INgbqf-xl07Ob-LgbsSe-hFsbo-L6cTce.VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { padding-right: 4px; }

.HB1eCd-MqDS2b-uoC0bf #replaceImageMenu .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { display: none; }

.HB1eCd-MqDS2b-uoC0bf #docs-align-palette { background: rgb(237, 242, 250); padding: 0px 4px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe .HB1eCd-Bz112c, .HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-LgbsSe .HB1eCd-Bz112c { height: 20px; margin-bottom: 0px; width: 20px; }

.HB1eCd-MqDS2b-uoC0bf .INgbqf-cjo6sd-Bz112c.HB1eCd-Bz112c { margin-bottom: -4px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m #docs-side-toolbar { margin-right: 12px; }

.HB1eCd-MqDS2b-uoC0bf #lineEndMenuButton .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed, .HB1eCd-MqDS2b-uoC0bf #lineStartMenuButton .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { margin-top: 0px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-hgDUwe.VIpgJd-TzA9Ye-eEGnhe { border-color: rgb(199, 199, 199); margin: 10px 3px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-INgbqf-z5C9Gb-LgbsSe-SmKAyb-Q4BLdf .HB1eCd-Bz112c { margin-left: 1px; }

.HB1eCd-MqDS2b-uoC0bf .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie + .VIpgJd-INgbqf-ornU0b-LgbsSe.VIpgJd-INgbqf-LgbsSe-barxie { border-radius: 4px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-INgbqf-nJjxad-Dd6Aae .VIpgJd-INgbqf-yiAvpe-LgbsSe-SmKAyb-Q4BLdf { margin: 0px 4px 0px 3px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-INgbqf-nJjxad-Dd6Aae .VIpgJd-INgbqf-yiAvpe-LgbsSe-YPqjbf { height: 28px !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed + .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd.HB1eCd-UMrnmb-hFsbo { padding: 0px 2px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .HB1eCd-k77Iif-IKhaXe .HB1eCd-UMrnmb-hFsbo.VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { margin: 1px -3px 0px -5px; }

.HB1eCd-MqDS2b-uoC0bf #headingStyleSelect .HB1eCd-UMrnmb-hFsbo, .HB1eCd-MqDS2b-uoC0bf #docs-font-family .HB1eCd-UMrnmb-hFsbo { margin: 0px 4px 0px 5px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { margin-left: 8px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-fmcmS-LgbsSe, .HB1eCd-MqDS2b-uoC0bf #docs-font-family .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { font-size: 14px; }

.HB1eCd-MqDS2b-uoC0bf #headingStyleSelect .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { font-size: 14px; width: 80px; }

.HB1eCd-MqDS2b-uoC0bf #docs-font-family .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { width: 55px; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-INgbqf-nJjxad-Dd6Aae .VIpgJd-INgbqf-yiAvpe-LgbsSe-cHYyed { width: 52px !important; }

.HB1eCd-MqDS2b-uoC0bf .HB1eCd-k77Iif-IKhaXe .HB1eCd-INgbqf-fmcmS-LgbsSe .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf { padding: 0px 8px; }

.HB1eCd-uWtm3-GMvhG-ORHb-Q3DXx-i8xkGf, .HB1eCd-uWtm3-GMvhG-ORHb-haAclf { align-items: center; display: flex; height: 40px; outline: none; overflow: hidden; width: 100%; }

.HB1eCd-uWtm3-GMvhG-ORHb-r4nke { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 15px; font-weight: 500; letter-spacing: 0.1px; margin: 0px 0px 0px 16px; }

.HB1eCd-uWtm3-GMvhG-ORHb-Ne3sFf { -webkit-box-flex: 1; flex-grow: 1; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; letter-spacing: 0.2px; margin: 0px 16px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.HB1eCd-uWtm3-GMvhG-ORHb-Bz112c { margin: 0px 0px 0px 16px; }

.HB1eCd-uWtm3-GMvhG-ORHb-c6xFrd { align-items: center; display: flex; }

.HB1eCd-uWtm3-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe { align-self: center; background-color: inherit; border: 1px inset transparent; border-radius: 100px; color: rgb(32, 33, 36); display: flex; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; line-height: 30px; outline: transparent solid 1px; padding: 0px 1px; text-transform: none; }

.HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe-haAclf .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe { border: 1px inset rgb(138, 180, 248); outline: rgb(210, 227, 252) solid 1px; border-radius: 4px; padding: 0px 1px; }

.HB1eCd-uWtm3-yJkfm-TZk80d-GMvhG-ORHb-haAclf, .HB1eCd-uWtm3-yJkfm-TZk80d-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-Q3DXx-i8xkGf { background-color: rgb(251, 188, 4); }

.HB1eCd-uWtm3-m9bMae-eKpHRd-QIk5de-GMvhG-ORHb-haAclf, .HB1eCd-uWtm3-m9bMae-eKpHRd-QIk5de-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-Q3DXx-i8xkGf { background-color: rgb(254, 247, 224); }

.HB1eCd-uWtm3-GMvhG-ORHb-JLm1tf-L7w45e-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc { box-shadow: rgb(32, 33, 36) 0px 0px 0px 1px; }

.HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc { border-radius: 100px; padding: 0px 24px; margin-top: 1px; margin-bottom: 1px; }

.HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc:hover { background-color: rgba(0, 0, 0, 0.12); }

.HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe-haAclf .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { background-color: transparent; }

.HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe-haAclf .HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e, .HB1eCd-uWtm3-GMvhG-ORHb-JIbuQc-LgbsSe-haAclf .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { line-height: 30px; border-radius: 100px; border: 1px inset transparent; outline: transparent solid 1px; padding: 0px 1px; }

.HB1eCd-uWtm3-yJkfm-TZk80d-oKM7Re-L7w45e-GMvhG-ORHb-haAclf, .HB1eCd-uWtm3-yJkfm-TZk80d-oKM7Re-L7w45e-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-Q3DXx-i8xkGf { background-color: rgb(179, 38, 30); color: rgb(255, 255, 255); }

.HB1eCd-uWtm3-yJkfm-TZk80d-oKM7Re-L7w45e-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JLm1tf-L7w45e-LgbsSe-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JLm1tf-L7w45e-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc, .HB1eCd-uWtm3-yJkfm-TZk80d-oKM7Re-L7w45e-GMvhG-ORHb-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JLm1tf-L7w45e-LgbsSe-haAclf .HB1eCd-uWtm3-GMvhG-ORHb-JLm1tf-L7w45e-LgbsSe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e .HB1eCd-HzV7m-LgbsSe-bN97Pc { color: rgb(255, 255, 255); box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px; }

#docs-omnibox-toolbar.nKilkd-LQLjdd-QbdDtf-L6cTce { display: none; }

#docs-omnibox-toolbar.nKilkd-LQLjdd { width: 100px; }

.HB1eCd-QbdDtf-YPqjbf.nKilkd-LQLjdd-INgbqf-QbdDtf { min-width: 98px; }

#docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-h0T7hb { position: fixed; width: 100px; }

#docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-h0T7hb .ztA2jd-oKdM2c .VIpgJd-j7LFlb { padding: 10px 15px 10px 35px; }

#docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-h0T7hb:focus-within { width: 350px; z-index: 1003; }

#docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd.nKilkd-LQLjdd-INgbqf-QbdDtf { padding-left: 35px; }

.HB1eCd-QbdDtf-h0T7hb .HB1eCd-QbdDtf-AaTFfe-clz4Ic { padding: 0.5em 0px; }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-auswjd .HB1eCd-QbdDtf-AaTFfe-clz4Ic { background-color: rgb(255, 255, 255); }

.HB1eCd-QbdDtf-h0T7hb .HB1eCd-QbdDtf-AaTFfe-clz4Ic .clz4Ic { margin: 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-YPqjbf:focus-within { border-radius: 8px 8px 0px 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd { padding: 0px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-Bz112c { margin: 4px 8px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-oKdM2c-Bz112c { margin: 1px 5px; }

.HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar .HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd[aria-expanded="true"].nKilkd-LQLjdd-INgbqf-QbdDtf { padding-left: 35px; }

.HB1eCd-MqDS2b-uoC0bf .nKilkd-LQLjdd-G0jgYd-LIIi-haAclf { gap: 1ch; display: flex; font-weight: 400; justify-content: center; }

.HB1eCd-MqDS2b-uoC0bf .nKilkd-LQLjdd-G0jgYd-LIIi-RmniWd-brjg8b { font-weight: 500; }

@media screen and (max-width: 1600px) {
  .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-YPqjbf { background-color: rgb(237, 242, 250); border-radius: 4px; }
  .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-YPqjbf { background-color: rgb(243, 246, 252); }
  .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-YPqjbf:hover { background-color: rgba(68, 71, 70, 0.08); cursor: pointer; padding-right: 0px; }
  .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-YPqjbf:focus-within { background: white; cursor: auto; }
  .HB1eCd-MqDS2b-uoC0bf .HB1eCd-QbdDtf-YPqjbf.nKilkd-LQLjdd-INgbqf-QbdDtf { min-width: 35px; }
  .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd, .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-h0T7hb { width: 35px; }
  .HB1eCd-MqDS2b-uoC0bf #docs-omnibox-toolbar.nKilkd-LQLjdd .HB1eCd-QbdDtf-h0T7hb:focus-within { width: 350px; }
}

#docs-meet-in-editors-entrypointbutton { background: rgb(255, 255, 255); border-radius: 33px; box-sizing: border-box; cursor: pointer; height: 36px; margin-right: 12px; width: 54px; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { cursor: default; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { box-shadow: none; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { background: rgb(241, 243, 244); border-color: rgb(241, 243, 244); }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background: rgb(232, 240, 254); border-color: rgb(232, 240, 254); }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-Bz112c { height: 24px; width: 24px; margin: 5px 4px 0px; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd .HB1eCd-Bz112c { margin-left: 8px; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c { background-color: rgb(26, 115, 232); border-radius: 100px; content: ""; height: 16px; margin: 4px auto 0px; position: initial; width: 4px; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c::before { background-color: rgb(26, 115, 232); border-radius: 100px; content: ""; display: inline-block; height: 8px; left: 4px; position: absolute; top: 8px; width: 4px; }

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c::after { background-color: rgb(26, 115, 232); border-radius: 100px; content: ""; display: inline-block; height: 8px; left: 16px; position: absolute; top: 8px; width: 4px; }

@media (forced-colors: active) {
  #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c, #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c::before, #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd-Bz112c::after { background-color: buttontext; }
}

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(26, 115, 232) transparent; right: 6px; top: 15px; }

@media (forced-colors: active) {
  #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: canvastext canvas; }
  @supports (forced-color-adjust: none) {
  #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { forced-color-adjust: none; border-color: canvastext transparent; }
}
}

#docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(32, 33, 36) transparent; }

#docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border-color: rgb(220, 220, 220); }

#docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { display: none; }

#docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { opacity: 1; }

.HB1eCd-B8pEb-bEDTcc-HivRGb-xl07Ob { background: rgb(255, 255, 255); border-radius: 8px; border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; padding: 0px; width: 330px; }

#docs-meet-in-editors-loading.L6cTce { display: none; }

#docs-meet-in-editors-loading { height: 270px; display: flex; align-items: center; justify-content: center; }

#docs-meet-in-editors-loading .HB1eCd-aZ2wEe { align-items: center; display: flex; overflow: visible; }

#docs-meet-in-editors-loading .HB1eCd-vyDMJf-aZ2wEe { top: auto; }

#docs-meet-in-editors-error { color: rgb(95, 99, 104); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; line-height: 18px; padding: 16px; text-align: center; }

#docs-meet-in-editors-error > img { display: block; margin-left: auto; margin-right: auto; }

#docs-meet-in-editors-error > div { margin: 22px 34px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton { align-items: center; background: none; border: 1px solid transparent; display: flex; height: 40px; margin-right: 8px; padding-bottom: 2px; width: 68px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { width: 56px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { padding: 0px 0px 2px 2px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { padding-left: 5px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background: rgb(232, 235, 238); }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd { background: rgb(225, 227, 230); }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border-color: transparent; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { background: rgba(11, 87, 208, 0.08); }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background: rgba(11, 87, 208, 0.12); }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-aTv5jf-F75qrd .HB1eCd-Bz112c { margin-left: 3px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(68, 71, 70) transparent; right: 14px; top: 17px; }

.HB1eCd-MqDS2b-uoC0bf #docs-meet-in-editors-entrypointbutton.HB1eCd-B8pEb-bEDTcc-HivRGb-auswjd-F75qrd.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(11, 87, 208) transparent; }

#docs-omnibox-toolbar .HB1eCd-QbdDtf-h0T7hb { margin-right: 4px; }

.HB1eCd-QbdDtf-h0T7hb { margin-top: 4px; }

.HB1eCd-QbdDtf-YPqjbf { box-sizing: border-box; width: 100%; min-width: 289px; }

.HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; letter-spacing: 0.2px; line-height: 36px; background-color: rgb(241, 243, 244); border: 1px solid transparent; border-radius: 8px; box-shadow: none; color: rgb(32, 33, 36); height: 36px; padding: 1px 7px; }

.HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd::placeholder { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; letter-spacing: 0.2px; line-height: 36px; color: rgb(95, 99, 104); }

#docs-omnibox-toolbar .HB1eCd-Bz112c { margin: 3px; }

.HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd:focus { background-color: rgb(255, 255, 255); border: 1px solid transparent; box-shadow: rgba(32, 33, 36, 0.28) 0px 1px 6px; padding: 1px 7px; }

.HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd:active { background-color: rgb(255, 255, 255); border: 1px solid transparent; box-shadow: rgba(32, 33, 36, 0.28) 0px 1px 6px; padding: 1px 7px; }

.HB1eCd-QbdDtf-YPqjbf.tk3N6e-y4JFTd:focus[aria-expanded="true"] { border-color: transparent transparent rgb(232, 234, 237); border-style: solid; border-width: 1px; border-radius: 8px 8px 0px 0px; padding: 1px 7px; }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-SUR3Rd { background-color: rgb(255, 255, 255); border-color: transparent; border-radius: 0px 0px 8px 8px; border-style: solid; border-width: 0px 1px 1px; box-shadow: rgba(32, 33, 36, 0.28) 0px 4px 6px; outline: none medium; padding: 6px 0px; position: fixed; width: auto; z-index: 1003; }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-oKdM2c { padding: 0px; }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-oKdM2c .VIpgJd-j7LFlb { padding: calc(0.4em + 5px) calc(0.4em + 10px) calc(0.4em + 5px) calc(0.4em + 30px); }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-AHUcCb { font-weight: 500; }

.HB1eCd-QbdDtf-h0T7hb .ztA2jd-auswjd { background-color: rgb(241, 243, 244); }

.HB1eCd-QbdDtf-h0T7hb .HB1eCd-Bz112c { cursor: pointer; margin: 3px 3px 3px 5px; pointer-events: none; position: absolute; }

[class*="docs-hc"] .HB1eCd-QbdDtf-h0T7hb .ztA2jd-auswjd .VIpgJd-j7LFlb { border-color: transparent; border-style: dotted; border-width: 1px 0px; padding-top: 5px; padding-bottom: 5px; }

[class*="docs-hc"] .HB1eCd-PtzLtb.VIpgJd-j7LFlb .ztA2jd-oKdM2c .VIpgJd-j7LFlb .VIpgJd-j7LFlb-Bz112c { margin-top: 7px; }

[class*="docs-hc"] .HB1eCd-PtzLtb.VIpgJd-j7LFlb .ztA2jd-oKdM2c.ztA2jd-auswjd .VIpgJd-j7LFlb-Bz112c { margin-top: 6px; }

.HB1eCd-QbdDtf-oKdM2c-bN97Pc { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-QbdDtf-tlSJBe.VIpgJd-xl07Ob-BvBYQ .HB1eCd-PtzLtb.VIpgJd-j7LFlb { padding-left: 16px; }

.HB1eCd-QbdDtf-tlSJBe .HB1eCd-PtzLtb.VIpgJd-j7LFlb.VIpgJd-j7LFlb-sn54Q { background-color: rgb(255, 255, 255); border-color: rgb(255, 255, 255); }

.HB1eCd-QbdDtf-tlSJBe .HB1eCd-PtzLtb { outline: none; }

.HB1eCd-QbdDtf-N7Eqid-hSRGPd { color: rgb(66, 133, 244); font-size: 12px; padding-left: 260px; padding-right: 8px; padding-top: 1px; text-decoration: underline; user-select: none; }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe { background: rgb(255, 255, 255); box-sizing: border-box; border-radius: 33px; cursor: pointer; height: 30px; margin-right: 12px; min-width: 54px; width: 78px; }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { cursor: default; }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd, .HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { box-shadow: none; }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { background: rgb(241, 243, 244); border-color: rgb(95, 99, 104); }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .HB1eCd-Bz112c { margin: 6px 4px; }

.HB1eCd-bOjP2c-u014N-H6j5tf-rtUoue-Btuy5e { align-items: center; align-self: center; background-color: rgb(241, 243, 244); border-radius: 9px; box-sizing: border-box; display: flex; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 500; height: 18px; justify-content: center; min-width: 18px; padding: 0px 5px; }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe .HB1eCd-bOjP2c-u014N-H6j5tf-rtUoue-Btuy5e, .HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .HB1eCd-bOjP2c-u014N-H6j5tf-rtUoue-Btuy5e { background: rgb(218, 220, 224); }

.HB1eCd-bOjP2c-u014N-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { display: flex; height: 30px; }

.HB1eCd-bOjP2c-u014N-fbvM8b-V67aGc { display: flex; align-self: center; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 500; justify-content: center; margin-right: 2px; }

.eCwPFe-N7Eqid-gbaOCd-zUJ9re-wvGCSb-h0T7hb-oKdM2c { box-sizing: border-box; padding: 8px 4px; overflow-wrap: break-word; }

.IyROMc-JIbuQc-mJSDk-Bz112c { direction: ltr; text-align: left; overflow: hidden; position: relative; vertical-align: middle; }

.IyROMc-JIbuQc-mJSDk-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/shortcut_sprite1.png"); }

.IyROMc-JIbuQc-mJSDk-RJLb9c { height: 95px; position: absolute; width: 21px; }

.IyROMc-JIbuQc-mJSDk-a4fUwd { left: 0px; top: -63px; }

.IyROMc-JIbuQc-mJSDk-a4fUwd-HLvlvd { left: 0px; top: -21px; }

.IyROMc-JIbuQc-mJSDk-TvD9Pc-PvhD9 { left: 0px; top: -84px; }

.IyROMc-JIbuQc-mJSDk-G0jgYd { left: 0px; top: -42px; }

.IyROMc-JIbuQc-mJSDk-G0jgYd-HLvlvd { left: 0px; top: 0px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf { -webkit-box-align: center; align-items: center; background: none; display: flex; height: 21px; outline: 0px; position: relative; width: 35px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-PFprWc { transition-duration: 0.28s; transition-property: all; transition-timing-function: cubic-bezier(0.4, 0, 0.2, 1); left: 0px; right: inherit; top: 0px; will-change: background-color; background-color: rgb(241, 241, 241); border-radius: 100%; box-shadow: rgba(0, 0, 0, 0.12) 0px 0px 2px, rgba(0, 0, 0, 0.24) 0px 2px 4px; height: 20px; width: 20px; position: absolute; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-barxie .IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-PFprWc { left: inherit; right: 0px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-OWB6Me { cursor: not-allowed; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-u014N { background-color: rgb(0, 0, 0); border-radius: 7px; height: 14px; opacity: 0.26; width: 35px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-barxie .IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-u014N { opacity: 0.5; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-u014N, .IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-PFprWc { border: 1px solid transparent; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-XpnDCe { outline: transparent solid 1px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-XpnDCe .IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-PFprWc { box-shadow: rgba(0, 0, 0, 0.14) 0px 0px 4px, rgba(0, 0, 0, 0.28) 0px 4px 8px; }

.IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-haAclf-ZmdkE .IyROMc-vWsuo-HzV7m-nKQ6qf-ornU0b-PFprWc { box-shadow: rgba(0, 0, 0, 0.16) 0px 0px 6px, rgba(0, 0, 0, 0.32) 0px 6px 12px; }

.ztA2jd-SUR3Rd { font: 13px Arial, sans-serif; position: absolute; background: rgb(255, 255, 255); border: 1px solid rgb(102, 102, 102); box-shadow: rgba(102, 102, 102, 0.4) 2px 2px 2px; width: 300px; }

.ztA2jd-oKdM2c { cursor: pointer; padding: 0.4em; }

.ztA2jd-AHUcCb { font-weight: bold; }

.ztA2jd-auswjd { background-color: rgb(178, 180, 191); }

.tk3N6e-LgbsSe { border-radius: 2px; cursor: default; font-size: 11px; font-weight: bold; text-align: center; white-space: nowrap; margin-right: 16px; height: 27px; line-height: 27px; min-width: 54px; outline: 0px; padding: 0px 8px; }

.tk3N6e-LgbsSe-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; }

.tk3N6e-LgbsSe-gk6SMd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.tk3N6e-LgbsSe .tk3N6e-LgbsSe-RJLb9c { margin-top: -3px; vertical-align: middle; }

.tk3N6e-LgbsSe-V67aGc { margin-left: 5px; }

.tk3N6e-LgbsSe-roVxwc { min-width: 34px; padding: 0px; }

.tk3N6e-LgbsSe-vhaaFf-LK5yu, .tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 1; }

.tk3N6e-LgbsSe-vhaaFf-LK5yu.tk3N6e-LgbsSe-OWB6Me { z-index: 0; }

.tk3N6e-LgbsSe-barxie.tk3N6e-LgbsSe-vhaaFf-LK5yu, .tk3N6e-LgbsSe-barxie.tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 2; }

.tk3N6e-LgbsSe-vhaaFf-LK5yu:focus, .tk3N6e-LgbsSe-vhaaFf-qwU8Me:focus, .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-vhaaFf-LK5yu, .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 3; }

.tk3N6e-LgbsSe-vhaaFf-LK5yu { margin-left: -1px; border-bottom-left-radius: 0px; border-top-left-radius: 0px; }

.tk3N6e-LgbsSe-vhaaFf-qwU8Me { margin-right: 0px; border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.tk3N6e-LgbsSe.tk3N6e-LgbsSe-OWB6Me:active { box-shadow: none; }

.tk3N6e-LgbsSe-JIbuQc { box-shadow: none; background-color: rgb(77, 144, 254); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(71, 135, 237)); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(53, 122, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); border: 1px solid rgb(47, 91, 183); }

.tk3N6e-LgbsSe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-JbbQac-i5vt6e { box-shadow: none; outline: none; }

.tk3N6e-LgbsSe-JIbuQc:active { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; background: rgb(53, 122, 232); border: 1px solid rgb(47, 91, 183); }

.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(77, 144, 254); opacity: 0.5; }

.tk3N6e-LgbsSe-haDnnc { box-shadow: none; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); color: rgb(68, 68, 68); border: 1px solid rgba(0, 0, 0, 0.1); }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-ZmdkE, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-haDnnc:active, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-ZmdkE:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background: rgb(248, 248, 248); }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-gk6SMd, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-gk6SMd { background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-barxie, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-barxie { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-haDnnc:focus { border: 1px solid rgb(77, 144, 254); outline: none; }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid rgb(220, 220, 220); outline: none; }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.tk3N6e-LgbsSe-haDnnc .tk3N6e-LgbsSe-RJLb9c { opacity: 0.55; }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-barxie .tk3N6e-LgbsSe-RJLb9c, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-gk6SMd .tk3N6e-LgbsSe-RJLb9c, .tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-ZmdkE .tk3N6e-LgbsSe-RJLb9c { opacity: 0.9; }

.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me .tk3N6e-LgbsSe-RJLb9c { opacity: 0.333; }

.tk3N6e-LgbsSe-zTETae { box-shadow: none; background-color: rgb(61, 148, 0); background-image: -webkit-linear-gradient(top, rgb(61, 148, 0), rgb(57, 138, 0)); border: 1px solid rgb(41, 105, 29); color: rgb(255, 255, 255); text-shadow: rgba(0, 0, 0, 0.1) 0px 1px; }

.tk3N6e-LgbsSe-zTETae.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(54, 130, 0); background-image: -webkit-linear-gradient(top, rgb(61, 148, 0), rgb(54, 130, 0)); border: 1px solid rgb(45, 98, 0); text-shadow: rgba(0, 0, 0, 0.3) 0px 1px; }

.tk3N6e-LgbsSe-zTETae:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.tk3N6e-LgbsSe-zTETae.tk3N6e-LgbsSe-JbbQac-i5vt6e { box-shadow: none; outline: none; }

.tk3N6e-LgbsSe-zTETae:active { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; background: rgb(54, 130, 0); border: 1px solid rgb(45, 98, 0); }

.tk3N6e-LgbsSe-zTETae.tk3N6e-LgbsSe-OWB6Me { background: rgb(61, 148, 0); opacity: 0.5; }

.tk3N6e-LgbsSe-Kb3HCc { border-radius: 0px; border: 1px solid transparent; font-size: 13px; font-weight: normal; height: 21px; line-height: 21px; margin-right: 1px; min-width: 0px; padding: 0px; }

.tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-ZmdkE, .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-gk6SMd, .tk3N6e-LgbsSe-Kb3HCc:focus, .tk3N6e-LgbsSe-Kb3HCc:active { box-shadow: none; }

.tk3N6e-LgbsSe-Kb3HCc .tk3N6e-LgbsSe-RJLb9c { height: 21px; opacity: 0.55; width: 21px; }

.tk3N6e-LgbsSe-Kb3HCc .tk3N6e-LgbsSe-V67aGc { display: inline-block; margin: 0px; padding: 0px 1px; }

.tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-gk6SMd .tk3N6e-LgbsSe-RJLb9c, .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-ZmdkE .tk3N6e-LgbsSe-RJLb9c { opacity: 0.9; }

.tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-OWB6Me .tk3N6e-LgbsSe-RJLb9c { opacity: 0.333; }

.tk3N6e-LgbsSe-Kb3HCc:focus { border: 1px solid rgb(77, 144, 254); }

.tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid transparent; }

.tk3N6e-LgbsSe-yolsp { background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); height: 17px; line-height: 17px; min-width: 22px; text-shadow: rgba(0, 0, 0, 0.1) 0px 1px; }

.tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-ZmdkE, .tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); text-shadow: rgba(0, 0, 0, 0.3) 0px 1px; }

.tk3N6e-LgbsSe-yolsp:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-barxie, .tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-barxie { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(224, 224, 224); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-yolsp:focus { border: 1px solid rgb(77, 144, 254); }

.tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid rgb(220, 220, 220); }

.tk3N6e-LgbsSe-yolsp.tk3N6e-LgbsSe-OWB6Me { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.tk3N6e-LgbsSe-ssJRIf { box-shadow: none; background-color: rgb(209, 72, 54); background-image: -webkit-linear-gradient(top, rgb(221, 75, 57), rgb(209, 72, 54)); border: 1px solid transparent; color: rgb(255, 255, 255); text-shadow: rgba(0, 0, 0, 0.1) 0px 1px; text-transform: uppercase; }

.tk3N6e-LgbsSe-ssJRIf.tk3N6e-LgbsSe-ZmdkE { box-shadow: rgba(0, 0, 0, 0.2) 0px 1px 1px; background-color: rgb(197, 55, 39); background-image: -webkit-linear-gradient(top, rgb(221, 75, 57), rgb(197, 55, 39)); border-width: 1px; border-style: solid; border-color: rgb(176, 40, 26) rgb(176, 40, 26) rgb(175, 48, 31); border-image: initial; }

.tk3N6e-LgbsSe-ssJRIf:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.tk3N6e-LgbsSe-ssJRIf.tk3N6e-LgbsSe-JbbQac-i5vt6e { box-shadow: none; outline: none; }

.tk3N6e-LgbsSe-ssJRIf:active { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; background-color: rgb(176, 40, 26); background-image: -webkit-linear-gradient(top, rgb(221, 75, 57), rgb(176, 40, 26)); border: 1px solid rgb(153, 42, 27); }

.tk3N6e-LgbsSe-ssJRIf.tk3N6e-LgbsSe-OWB6Me { background: rgb(209, 72, 54); opacity: 0.5; }

.tk3N6e-LR6Drb { border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px 0px inset; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border: 1px solid rgb(204, 204, 204); color: rgb(102, 102, 102); font-weight: bold; height: 27px; line-height: 27px; margin-right: 16px; outline: none; overflow: hidden; padding: 0px; position: relative; width: 94px; }

.tk3N6e-LR6Drb-IT5dJd, .tk3N6e-LR6Drb-Xhs9z, .tk3N6e-LR6Drb-PFprWc { display: inline-block; text-align: center; text-transform: uppercase; width: 47px; }

.tk3N6e-LR6Drb-IT5dJd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px 0px inset; background-color: rgb(57, 139, 242); background-image: -webkit-linear-gradient(top, rgb(59, 147, 255), rgb(54, 137, 238)); color: rgb(255, 255, 255); height: 27px; }

.tk3N6e-LR6Drb-Xhs9z { border-radius: 2px 2px 0px 0px; }

.tk3N6e-LR6Drb-PFprWc { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px 0px; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); transition: all 0.13s ease-out 0s; border: 1px solid rgb(204, 204, 204); display: block; height: 27px; left: -1px; position: absolute; top: -1px; }

.tk3N6e-LR6Drb-PFprWc::after { content: ""; background-position: 0px 0px, 0px 2px, 0px 4px, 0px 6px, 0px 8px; background-repeat: repeat-x; background-size: 2px 1px; display: block; height: 9px; left: 15px; position: absolute; top: 9px; width: 17px; }

.tk3N6e-LR6Drb.tk3N6e-LR6Drb-barxie .tk3N6e-LR6Drb-PFprWc { left: 47px; }

.tk3N6e-LR6Drb:focus { border: 1px solid rgb(77, 144, 254); }

.tk3N6e-LR6Drb.tk3N6e-LR6Drb-kyhDef { border: 1px solid rgb(204, 204, 204); }

.tk3N6e-LgbsSe-n2to0e { box-shadow: none; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); color: rgb(68, 68, 68); border: 1px solid rgba(0, 0, 0, 0.1); }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-n2to0e:active, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background: rgb(248, 248, 248); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-gk6SMd, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-gk6SMd { background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-barxie, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-barxie { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.tk3N6e-LgbsSe-n2to0e:focus { border: 1px solid rgb(77, 144, 254); outline: none; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid rgba(0, 0, 0, 0.1); outline: none; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.tk3N6e-LgbsSe-n2to0e .tk3N6e-LgbsSe-RJLb9c { opacity: 0.55; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-barxie .tk3N6e-LgbsSe-RJLb9c, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-gk6SMd .tk3N6e-LgbsSe-RJLb9c, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE .tk3N6e-LgbsSe-RJLb9c { opacity: 0.9; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me .tk3N6e-LgbsSe-RJLb9c { opacity: 0.333; }

.VIpgJd-TUo6Hb, .XKSfm-Sx9Kwc { box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; background: padding-box rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.333); outline: 0px; position: absolute; }

.VIpgJd-TUo6Hb-xJ5Hnf, .XKSfm-Sx9Kwc-xJ5Hnf { background: rgb(255, 255, 255); left: 0px; position: absolute; top: 0px; }

div.VIpgJd-TUo6Hb-xJ5Hnf, div.XKSfm-Sx9Kwc-xJ5Hnf { opacity: 0.75; }

.XKSfm-Sx9Kwc { color: rgb(0, 0, 0); padding: 30px 42px; }

.XKSfm-Sx9Kwc-r4nke { background-color: rgb(255, 255, 255); color: rgb(0, 0, 0); cursor: default; font-size: 16px; font-weight: normal; line-height: 24px; margin: 0px 0px 16px; }

.XKSfm-Sx9Kwc-r4nke-TvD9Pc { height: 11px; opacity: 0.7; padding: 17px; position: absolute; right: 0px; top: 0px; width: 11px; }

.XKSfm-Sx9Kwc-r4nke-TvD9Pc::after { content: ""; background: url("//ssl.gstatic.com/ui/v1/dialog/close-x.png"); position: absolute; height: 11px; width: 11px; right: 17px; }

.XKSfm-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.XKSfm-Sx9Kwc-bN97Pc { background-color: rgb(255, 255, 255); line-height: 1.4em; overflow-wrap: break-word; }

.XKSfm-Sx9Kwc-c6xFrd { margin-top: 16px; }

.XKSfm-Sx9Kwc-c6xFrd button { border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); cursor: default; font-family: inherit; font-size: 11px; font-weight: bold; height: 29px; line-height: 27px; margin: 0px 16px 0px 0px; min-width: 72px; outline: 0px; padding: 0px 8px; }

.XKSfm-Sx9Kwc-c6xFrd button:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.XKSfm-Sx9Kwc-c6xFrd button:active { background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.XKSfm-Sx9Kwc-c6xFrd button:focus { border: 1px solid rgb(77, 144, 254); }

.XKSfm-Sx9Kwc-c6xFrd button[disabled] { box-shadow: none; background: none rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc { background-color: rgb(77, 144, 254); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(71, 135, 237)); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover { background-color: rgb(53, 122, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); }

.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active { background-color: rgb(53, 122, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; }

.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled] { box-shadow: none; background: rgb(77, 144, 254); color: rgb(255, 255, 255); opacity: 0.5; }

.tk3N6e-O0r3Gd, .tk3N6e-McfNlf, .tk3N6e-ostUZ { width: 512px; }

.tk3N6e-y4JFTd { border-radius: 1px; border-width: 1px; border-style: solid; border-color: rgb(192, 192, 192) rgb(217, 217, 217) rgb(217, 217, 217); border-image: initial; font-size: 13px; height: 25px; padding: 1px 8px; }

.tk3N6e-y4JFTd:focus { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; border: 1px solid rgb(77, 144, 254); outline: none; }

.IyROMc-w3KqTd { top: 0px; z-index: 1002; color: rgb(33, 33, 33); font-family: roboto, arial, sans-serif; font-size: 13px; position: fixed; text-align: center; background: none 0px center repeat scroll rgb(250, 250, 250); overflow: hidden; box-shadow: rgba(255, 255, 255, 0.9) 0px 1px 0px inset, rgba(0, 0, 0, 0.03) 0px -1px 0px inset, rgba(0, 0, 0, 0.15) 0px 15px 10px, rgba(0, 0, 0, 0.3) 0px 8px 36px; border: 1px solid transparent; }

.IyROMc-w3KqTd input { font-family: roboto, arial, sans-serif; }

@media print {
  .IyROMc-w3KqTd { display: none; }
}

.IyROMc-w3KqTd-xJ5Hnf { display: none; left: 0px; top: 0px; position: absolute; }

.IyROMc-w3KqTd-haAclf { display: flex; flex-direction: column; box-sizing: border-box; padding: 16px 32px; width: 800px; height: 600px; }

.IyROMc-w3KqTd-tJHJj, .IyROMc-w3KqTd-bN97Pc { border-collapse: collapse; width: 100%; }

.IyROMc-w3KqTd-tJHJj { flex: 0 0 auto; border-bottom: 1px solid rgb(229, 229, 229); text-align: left; }

.IyROMc-w3KqTd-bN97Pc { font-size: 13px; outline-offset: -1px; }

.IyROMc-w3KqTd-tJHJj-PQbLGe { display: inline-block; vertical-align: middle; height: 48px; }

.IyROMc-w3KqTd-r4nke-haAclf { white-space: nowrap; text-align: left; }

.IyROMc-w3KqTd-Sx9Kwc-r4nke { font-size: 16px; color: rgb(33, 33, 33); display: inline-block; vertical-align: middle; }

.IyROMc-w3KqTd-YPqjbf { font-size: 13px; margin-left: 16px; margin-right: 0px; padding: 0px 5px; vertical-align: middle; border-right: none; width: 250px; height: 27px; box-sizing: border-box; }

.IyROMc-w3KqTd-YPqjbf-LgbsSe-RJLb9c { height: 21px; width: 21px; display: inline-block; }

.IyROMc-w3KqTd-YPqjbf-LgbsSe { box-sizing: border-box; cursor: pointer; display: inline-block; margin-left: 0px; vertical-align: middle; border-top-left-radius: 0px; border-bottom-left-radius: 0px; line-height: 25px; }

.IyROMc-w3KqTd-tCq0Eb-hSRGPd { font-size: 13px; cursor: pointer; text-decoration: underline; color: rgb(69, 129, 255); vertical-align: middle; display: block; padding: 16px 0px 13px; font-weight: bold; }

.IyROMc-w3KqTd-TvD9Pc { position: absolute; top: 0px; right: 0px; padding-right: 30px; padding-top: 30px; }

.IyROMc-w3KqTd-TvD9Pc svg { fill: rgb(95, 99, 104); }

.IyROMc-w3KqTd-TvD9Pc-DH6Rkf-m5SR9c-qnnXGd { padding-right: 18px; padding-top: 20px; }

.IyROMc-w3KqTd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc { cursor: pointer; position: static; padding: 0px; margin: 0px 0px 0px 32px; vertical-align: middle; }

.IyROMc-w3KqTd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc::after { background: none; display: none; }

.IyROMc-w3KqTd-G0jgYd-ORHb { flex: 0 0 auto; text-align: left; height: 48px; padding-top: 12px; box-sizing: border-box; }

.IyROMc-w3KqTd-G0jgYd-ORHb.IyROMc-w3KqTd-xFQqWe-G0jgYd { position: relative; left: 0px; right: 0px; text-align: center; top: 113px; height: 48px; }

.IyROMc-w3KqTd-S9gUrf-G0jgYd-LgbsSe { cursor: pointer; text-decoration: underline; position: relative; width: 21px; min-width: 21px; display: inline-block; margin-right: 8px; }

.IyROMc-w3KqTd-S9gUrf-G0jgYd-LgbsSe-Bz112c { height: 21px; width: 21px; }

.IyROMc-w3KqTd-G0jgYd-V67aGc { margin: 0px; position: relative; font-size: 15px; display: inline-block; vertical-align: middle; }

.IyROMc-w3KqTd-aVTXAb-haAclf { flex: 1 1 auto; overflow: auto; }

.IyROMc-w3KqTd-bN97Pc-tJHJj { height: 48px; padding-top: 25px; text-align: left; font-size: 13px; color: rgb(33, 33, 33); white-space: nowrap; margin: 0px; box-sizing: border-box; }

.IyROMc-w3KqTd-bN97Pc-tJHJj.IyROMc-w3KqTd-bN97Pc-tJHJj-r08add { height: 32px; padding-top: 8px; }

.IyROMc-w3KqTd-bN97Pc-PQbLGe { text-align: left; vertical-align: middle; padding-top: 0.15em; border-bottom: 1px solid rgb(236, 236, 236); height: 32px; white-space: nowrap; box-sizing: border-box; }

.IyROMc-w3KqTd-mJSDk-Dzid5 { color: rgb(117, 117, 117); }

.IyROMc-w3KqTd-mJSDk-tEE2Ac { font-weight: bold; }

.IyROMc-w3KqTd-ztA2jd-SUR3Rd { z-index: 1003; font-family: Arial, sans-serif; font-size: 13px; position: absolute; background: rgb(255, 255, 255); border: 1px solid rgb(102, 102, 102); box-shadow: rgba(102, 102, 102, 0.4) 2px 2px 2px; width: 250px; box-sizing: border-box; }

.IyROMc-w3KqTd-ztA2jd-oKdM2c { cursor: pointer; padding: 0.4em; }

.IyROMc-w3KqTd-ztA2jd-SUR3Rd .ztA2jd-auswjd { background-color: rgb(238, 238, 238); }

.auswjd-mzNpsf-Sx9Kwc-xvr5H { font-weight: 500; word-break: break-all; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { display: flex; }

.auswjd-mzNpsf-Sx9Kwc-KVuj8d-V1ur5d { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; line-height: 12px; padding: 8px; display: flex; align-items: center; }

.auswjd-mzNpsf-Sx9Kwc-YLEF4c { background-color: rgb(154, 160, 166); border-radius: 50%; object-fit: cover; height: 32px; width: 32px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd { margin-top: 32px; }

.XKSfm-Sx9Kwc.auswjd-mzNpsf-Sx9Kwc { display: table; max-width: 464px; table-layout: fixed; }

.ndfHFb-c4YZDc-K9a4Re { position: absolute; transition: bottom 0.218s ease-out 0s; inset: 0px; z-index: 0; }

.fFW7wc-L5Fo6c.fFW7wc-jJNx8e { box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; color: rgb(0, 0, 0); padding: 0px; position: absolute; z-index: 1002; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-OEVmcd-yHKmmc { background-color: rgb(241, 241, 241); }

.fFW7wc-L5Fo6c.fFW7wc-HLvlvd-Hn6s1b.fFW7wc-VWkKje .fFW7wc-jJNx8e-OEVmcd-yHKmmc { background-color: rgb(255, 255, 255); }

.fFW7wc-L5Fo6c.fFW7wc-jJNx8e.VIpgJd-xl07Ob { border-color: rgb(204, 204, 204); line-height: 0; max-height: none; overflow: visible; }

.fFW7wc-L5Fo6c.fFW7wc-jJNx8e-ma6Yeb { margin-top: 15px; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje.fFW7wc-jJNx8e-ma6Yeb { margin-top: 9px; }

.fFW7wc-L5Fo6c.fFW7wc-jJNx8e-cGMI2b { margin-top: -15px; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje.fFW7wc-jJNx8e-cGMI2b { margin-top: -9px; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc, .fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW { position: absolute; width: 32px; z-index: 0; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc { top: -15px; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc { top: -10px; width: 20px; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW { bottom: -16px; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-hgHJW { bottom: -10px; width: 20px; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-SmKAyb, .fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-VtOx3e { border: 16px solid; height: 0px; position: absolute; width: 0px; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-SmKAyb, .fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-VtOx3e { border: 10px solid; }

.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb { border-color: rgb(241, 241, 241) transparent; }

.fFW7wc-L5Fo6c.fFW7wc-HLvlvd-Hn6s1b.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb { border-color: rgb(255, 255, 255) transparent; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb { border-color: rgb(255, 255, 255) transparent; top: 1px; z-index: 1; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-SmKAyb { border-color: rgb(255, 255, 255) transparent; bottom: 1px; z-index: 1; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-VtOx3e { border-color: rgba(0, 0, 0, 0.2) transparent; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-VtOx3e { border-color: rgba(0, 0, 0, 0.2) transparent; bottom: 0px; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb, .fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-VtOx3e { border-top-width: 0px; }

.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-SmKAyb, .fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-VtOx3e { border-bottom-width: 0px; }

.ndfHFb-c4YZDc { color: rgb(255, 255, 255); font-family: arial, sans-serif; overflow: clip; opacity: 0; visibility: hidden; transition: opacity 0.1s cubic-bezier(0, 0, 0.2, 1) 0s, visibility 0s 0.1s; position: fixed; inset: 0px; z-index: 100; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb { font-family: "Google Sans", Roboto, arial, sans-serif; }

.ndfHFb-c4YZDc-TSZdd { opacity: 1; visibility: visible; transition-timing-function: cubic-bezier(0.4, 0, 1, 1); transition-delay: 0s, 0s; }

.ndfHFb-c4YZDc-bnBfGc { background-color: rgb(30, 30, 30); position: fixed; inset: 0px; opacity: 0.93; }

.ndfHFb-c4YZDc-JNEHMb { left: 0px; position: absolute; right: 0px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-bnBfGc { background-color: rgb(209, 209, 209); opacity: 1; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bnBfGc { background-color: rgba(0, 0, 0, 0.85); opacity: 1; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bnBfGc { background-color: rgba(31, 31, 31, 0.92); }

.ndfHFb-c4YZDc-qbOKL-OEVmcd { margin: 0px; height: 100%; width: 100%; overflow: hidden !important; }

.ndfHFb-c4YZDc-AHmuwe-Hr88gd-OWB6Me :focus { outline: none; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc { display: flex; flex-direction: column; align-items: flex-start; padding-bottom: 16px; outline: none; position: absolute; width: 384px; height: auto; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; border-radius: 8px; z-index: 102; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-bN97Pc { max-width: 100%; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); height: 100%; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 101; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-r4nke { margin: 0px auto; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -64px; width: 24px; height: 24px; margin: 18px auto 10px; transform: scale(1.3); }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1.375rem; font-weight: 400; letter-spacing: 0px; line-height: 1.75rem; color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-C7uZwb-bN97Pc { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; display: flex; height: 100px; flex-direction: column; margin: 16px 24px 20px; justify-content: space-around; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-hSRGPd { color: rgb(95, 99, 104); overflow: hidden; text-overflow: ellipsis; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-Ne3sFf { color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-KY1xSc-z5C9Gb { font-weight: 100; margin: 0px 5px; position: relative; top: -2px; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-c6xFrd { margin-left: auto; margin-right: 24px; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-ssJRIf-LgbsSe:hover, .ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-K4efff-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-ssJRIf-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; text-align: center; min-width: 70px; background: rgb(249, 171, 0); border-radius: 5px; font-size: 14px; padding: 8px 24px; border-style: none; outline: none; }

.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-K4efff-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; margin: 0px 16px; text-align: center; min-width: 70px; font-size: 14px; padding: 7px 0px; border-style: none; background: rgb(255, 255, 255); outline: none; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { color: rgba(255, 255, 255, 0.87); font-size: 11px; font-weight: bold; text-align: center; text-shadow: rgba(0, 0, 0, 0.8) 0px 1px 0px; vertical-align: middle; height: 27px; line-height: 27px; margin-right: 2px; min-width: 50px; padding: 10px 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { text-shadow: none; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { border-radius: 2px; height: 24px; line-height: 24px; margin: 0px; padding: 8px; min-width: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { border-radius: 100px; }

.ndfHFb-c4YZDc-AHmuwe-Hr88gd-qnnXGd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { border-color: rgb(87, 87, 87); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-AHmuwe-Hr88gd-qnnXGd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { background-color: rgba(196, 199, 197, 0.12); }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me { color: rgba(255, 255, 255, 0.47); text-shadow: none; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background-color: rgb(35, 35, 35); background-image: -webkit-linear-gradient(top, rgb(51, 51, 51), rgb(34, 34, 34)); }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgb(131, 131, 131); background-image: none; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.8) 0px 1px 6px inset; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-LgbsSe-auswjd { box-shadow: none; background-color: rgba(255, 255, 255, 0.35); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-LgbsSe-auswjd { background-color: rgba(196, 199, 197, 0.12); }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe { background-color: rgba(35, 35, 35, 0.6); border-bottom: 3px solid rgb(77, 144, 254); padding-bottom: 7px; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe { background-color: rgb(109, 110, 113); border-bottom-color: rgb(88, 89, 91); }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgb(131, 131, 131); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { transition: background-color 0.1s ease 0s, opacity 0.1s ease 0s; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe .ndfHFb-c4YZDc-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgba(255, 255, 255, 0.25); background-image: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgba(196, 199, 197, 0.08); }

.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe, .ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe { background-color: rgba(255, 255, 255, 0.1); border-bottom-color: rgb(193, 217, 255); }

.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd, .ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.4) 0px 1px 6px inset; }

.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE, .ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE, .ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe, .ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { background: rgb(96, 156, 253); outline: 0px; }

.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { background: rgb(31, 89, 192); }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd { display: inline-block; margin: 6px 0px; }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe { background-color: rgb(63, 118, 217); }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background: rgb(64, 127, 241); }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac.ndfHFb-c4YZDc-to915-LgbsSe { margin-right: 1px; min-width: 35px; width: 35px; padding: 4px 0px; margin-left: 5px; }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac .ndfHFb-c4YZDc-Bz112c { background-position: 0px 0px; width: 25px; height: 25px; padding: 3px 10px; margin-left: 4px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1528px; }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-V67aGc { font-size: 13px; text-transform: uppercase; text-shadow: none; color: white; display: inline-block; padding-left: 3px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-Wrql6b-gvZm2b-xl07Ob-LgbsSe { padding: 4px 10px; margin-right: 5px; }

.ndfHFb-c4YZDc-Wrql6b-gvZm2b-xl07Ob-LgbsSe .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo { margin-left: 5px; }

.ndfHFb-c4YZDc .ndfHFb-aZ2wEe { display: none; height: 100%; width: 100%; }

.ndfHFb-c4YZDc .ndfHFb-vyDMJf-aZ2wEe { height: 21px; margin-left: -10.5px; top: 0px; width: 21px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-vyDMJf-aZ2wEe { height: 24px; margin-left: -12px; width: 24px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb { display: inline-block; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb { z-index: 1; display: none; }

.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c { background-repeat: no-repeat; opacity: 0.87; margin-left: auto; margin-right: auto; margin-top: 3px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c { background-repeat: no-repeat; opacity: 0.87; margin-left: auto; margin-right: auto; height: 21px; }

.ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c { background-repeat: no-repeat; opacity: 0.87; margin-left: auto; margin-right: auto; margin-top: 3px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c, .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c, .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c { background-repeat: no-repeat; opacity: 0.87; margin-left: auto; margin-right: auto; margin-top: 2px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg") !important; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-spinner_dark.gif") !important; }

.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c { background-position: 0px -240px; }

.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c { background-position: 0px -600px; }

.ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c { background-position: 0px -400px; }

.ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c { background-position: 0px -1920px; }

.ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c { margin-top: 4px; width: 19px; }

.ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c { background-position: 0px -2360px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited) { margin-top: 2px; height: 24px; width: 24px; opacity: 1; background-image: none !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c .ndfHFb-aZ2wEe { display: block; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg") !important; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c { background-position: 0px -1816px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c { background-position: 0px -1448px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c { background-position: 0px -896px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c { background-position: 0px -1568px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c { background-position: 0px -448px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c { background-position: 0px -328px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c { background-position: 0px -2464px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c { opacity: 1; margin-top: 0px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c { opacity: 1; margin: 2.5px; width: 19px; height: 19px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited) { margin: 0px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-Sx9Kwc.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc { padding: 0px; }

.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-r4nke { border-bottom: 1px solid rgb(172, 172, 172); font-family: arial, sans-serif; padding: 15px 12px; }

.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde { background-color: rgb(243, 243, 243); height: 100%; position: relative; width: 100%; }

.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde .ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde-k4Qmrd { text-align: center; width: 100%; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-ge6pde-RJLb9c { background-image: url("//ssl.gstatic.com/ui/v1/activityindicator/loading_bg_f5.gif"); background-repeat: no-repeat; display: inline-block; height: 19px; position: relative; top: 3px; width: 19px; }

.ndfHFb-c4YZDc-y0R6E-DWWcKd-b3rLgd { display: inline-block; vertical-align: middle; }

.ndfHFb-c4YZDc-y0R6E-DWWcKd-Bz112c { display: inline-block; height: 12px; width: 12px; }

.ndfHFb-c4YZDc-y0R6E-DWWcKd-Ne3sFf { display: inline-block; padding-left: 16px; vertical-align: top; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-xJ5Hnf { background-color: rgb(32, 33, 36); left: 0px; position: absolute; top: 0px; z-index: 101; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc { background-color: rgb(255, 255, 255); border-radius: 8px; font-family: "Google Sans", Roboto, arial, sans-serif; padding: 20px; position: absolute; width: 450px; z-index: 102; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-c6xFrd { float: right; margin-top: 20px; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-LgbsSe { background: rgb(255, 255, 255); border-color: rgb(189, 193, 198); border-radius: 4px; border-style: solid; border-width: 1px; color: rgb(26, 115, 232); cursor: pointer; font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 2; margin-left: 5px; padding: 0px 20px; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-zTETae { background: rgb(26, 115, 232); color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-r4nke-fmcmS { font-size: 22px; }

.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-bN97Pc { color: rgb(95, 99, 104); font-size: 14px; margin: 10px 0px; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf { display: none; align-items: center; background: rgb(232, 240, 254); color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, arial, sans-serif; height: 48px; width: 100%; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf { background: rgb(124, 172, 248); }

.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf.ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce, .ndfHFb-c4YZDc-MqcBrc-ORHb-c6xFrd.ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce, .ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce { display: none; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-c6xFrd { align-items: center; display: flex; -webkit-box-flex: 1; flex-grow: 1; float: right; justify-content: flex-end; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-Bz112c { background-position: 0px -2544px; height: 24px; margin: 0px 16px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-Bz112c { background-position: 0px -3634px; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-Vkfede-Ne3sFf { margin-left: 16px; font-size: 14px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-Vkfede-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-MqcBrc-ORHb-jOfkMb { font-size: 16px; font-weight: 500; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-jOfkMb { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); }

.ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-Bz112c { background-position: 0px -1160px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-Bz112c { background-position: 0px -3570px; height: 20px; width: 24px; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-sM5MNb { margin: 0px 16px; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover, .ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe { margin: 0px 12px; text-align: center; min-width: 70px; background: rgb(26, 115, 232); border-radius: 5px; font-size: 14px; font-weight: 500; padding: 7px 0px; color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe { margin: 0px 12px; color: rgb(32, 33, 36); background: none; font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); }

.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover { background: rgb(43, 125, 233); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover { background: none; }

.ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe { margin: 0px 5px; text-align: center; min-width: 70px; color: rgb(26, 115, 232); font-size: 14px; font-weight: 500; padding: 7px 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe { margin: 0px 12px; color: rgb(32, 33, 36); background: none; font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); }

.ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover { background: rgb(248, 251, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover { background: none; }

.ndfHFb-c4YZDc-rovI0b { color: rgb(255, 255, 255); font-size: 13px; font-weight: normal; text-align: left; text-shadow: rgba(0, 0, 0, 0.1) 0px 2px 1px; white-space: nowrap; }

.ndfHFb-c4YZDc-rovI0b-r4nke { line-height: 30px; margin-bottom: 10px; text-align: center; }

.ndfHFb-c4YZDc-rovI0b-bN97Pc { overflow: hidden auto; border-top: 1px solid rgb(105, 104, 104); border-bottom: 1px solid rgb(105, 104, 104); min-height: 55px; }

.ndfHFb-c4YZDc-rovI0b-bN97Pc.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb { min-height: 0px !important; }

.ndfHFb-c4YZDc-rovI0b-LS81yb { padding-bottom: 10px; }

.ndfHFb-c4YZDc-rovI0b-LS81yb-Ud7fr { border-bottom: none; color: rgb(205, 205, 205); font-size: 13px; font-weight: normal; line-height: 25px; padding: 0px; }

.ndfHFb-c4YZDc-rovI0b-IyROMc-rymPhb { margin-left: 100px; }

.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b { cursor: pointer; display: block; padding: 6px 15px 6px 0px; border: none; }

.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b.ndfHFb-c4YZDc-w5vlXd { border: none; }

.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b:hover { background-color: rgb(68, 68, 68); border-color: rgb(68, 68, 68); border-style: dotted; border-width: 1px 0px; padding: 5px 15px 5px 0px; }

.ndfHFb-c4YZDc-rovI0b-ljLd3-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b { font-weight: bold; }

.ndfHFb-c4YZDc-rovI0b-UEIKff-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b, .ndfHFb-c4YZDc-rovI0b-MVH0Ye-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b { font-weight: normal; }

.ndfHFb-c4YZDc-rovI0b-DWWcKd-Bz112c { display: inline-block; height: 16px; margin-left: 5px; vertical-align: middle; width: 16px; }

.ndfHFb-c4YZDc-rovI0b-DWWcKd-V1ur5d { display: inline-block; line-height: 16px; margin-left: 20px; }

.ndfHFb-c4YZDc-JqEhuc-s2gQvd { bottom: 0px; overflow: auto; position: absolute; }

.ndfHFb-c4YZDc-JqEhuc { background-color: rgb(255, 255, 255); border: 20px solid transparent; border-radius: 20px; color: rgb(0, 0, 0); font-size: 14px; position: absolute; overflow-wrap: break-word; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-JqEhuc { border-right: none; border-bottom: none; border-left: none; border-image: initial; border-radius: 0px; border-top: 10px solid transparent; box-shadow: none; }

.ndfHFb-c4YZDc-JqEhuc-bN97Pc, .ndfHFb-c4YZDc-JqEhuc-tJHJj { margin-left: 20px; margin-right: 20px; right: 0px; left: 0px; }

.ndfHFb-c4YZDc-JqEhuc-n5VRYe { background-image: linear-gradient(rgba(0, 0, 0, 0.2), transparent); height: 8px; left: 20px; position: absolute; right: 20px; z-index: 1; -webkit-mask-box-image-source: -webkit-linear-gradient(left, rgba(0, 0, 0, 0.1), rgba(0, 0, 0, 0.8), rgba(0, 0, 0, 0.8), rgba(0, 0, 0, 0.1)); -webkit-mask-box-image-slice: initial; -webkit-mask-box-image-width: initial; -webkit-mask-box-image-outset: initial; -webkit-mask-box-image-repeat: initial; }

.ndfHFb-c4YZDc-JqEhuc-r4nke { display: inline-block; font-size: 30px; margin-right: 10px; margin-left: 10px; max-width: 85%; opacity: 0.6; overflow: hidden; padding-bottom: 10px; text-overflow: ellipsis; vertical-align: middle; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-r4nke { line-height: 50px; padding-bottom: 0px; }

.ndfHFb-c4YZDc-JqEhuc-r4nke-tJHJj { border-bottom: 1px solid rgb(206, 206, 207); }

.ndfHFb-c4YZDc-JqEhuc-r4nke-oKdM2c { opacity: 0.6; font-size: 10px; display: block; overflow: hidden; white-space: nowrap; }

.ndfHFb-c4YZDc-JqEhuc-NnAfwf { display: inline-block; font-size: 16px; opacity: 0.6; vertical-align: middle; }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c, .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c { border-bottom: 1px solid rgb(206, 206, 207); display: block; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c.ndfHFb-c4YZDc-LgbsSe { display: block; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-tJHJj .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c { height: 50px; }

.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe, .ndfHFb-c4YZDc-JqEhuc-PlOyMe-Bz112c.ndfHFb-c4YZDc-LgbsSe, .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-JqEhuc-oKdM2c, .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c { cursor: pointer; }

.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-JqEhuc-oKdM2c, .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c, .ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe:hover, .ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe:active, .ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { background-color: rgb(221, 221, 221); }

.ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-oKdM2c, .ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-bMcfAe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-oKdM2c, .ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c, .ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-bMcfAe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c { background-color: rgb(232, 240, 254); color: rgb(24, 90, 188); }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c-Bz112c { background-size: contain; display: inline-block; height: 16px; width: 16px; margin-left: 10px; margin-right: 10px; position: relative; top: 3px; }

.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-Bz112c { background-size: contain; display: inline-block; height: 16px; width: 16px; margin-left: 3%; margin-right: 3%; position: relative; top: 10px; }

.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c { background-position: 0px -1840px; height: 21px; width: 21px; left: -5px; top: 8px; position: absolute; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c { background-position: 0px -1080px; }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c-V1ur5d { display: inline; line-height: 38px; }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb { float: left; }

.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d, .ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd, .ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe { display: inline-block; line-height: 38px; overflow: hidden; text-overflow: ellipsis; }

.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d { width: 50%; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d { font-size: 12px; }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd { width: 22%; opacity: 0.6; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd { font-size: 12px; opacity: 1; }

.ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe { width: 13%; opacity: 0.6; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe { font-size: 12px; opacity: 1; }

.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c::after { content: ""; display: table; clear: both; }

.ndfHFb-c4YZDc-kODWGd { position: absolute; }

.ndfHFb-c4YZDc-kODWGd-nK2kYb { user-select: none; border-radius: 5px; background-color: rgba(20, 20, 20, 0.8); position: absolute; height: 100%; width: 100%; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; }

.ndfHFb-c4YZDc-kODWGd-NziyQe-LgbsSe { position: absolute; top: 2px; left: 10px; right: auto; }

.ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c { height: 28px; width: 26px; }

.ndfHFb-c4YZDc-kODWGd-NziyQe-Bz112c { height: 28px; width: 26px; background-position: 0px -1120px; }

.ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c { background-position: 0px -120px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-NziyQe-Bz112c { background-position: 0px -3386px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c { background-position: 0px -2344px; }

.ndfHFb-c4YZDc-kODWGd-bVEB4e { border: 1px solid rgb(179, 179, 179); background-color: rgb(10, 10, 10); display: table-cell; pointer-events: auto; text-align: center; vertical-align: middle; }

.ndfHFb-c4YZDc-kODWGd-LgbsSe { border-radius: 0px; transition: all 0.218s ease 0s; background-color: rgb(243, 243, 243); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); font-weight: bold; font-size: 11px; height: 27px; line-height: 27px; margin: 6px; min-width: 54px; padding: 0px 8px; text-align: center; }

.ndfHFb-c4YZDc-kODWGd-LgbsSe:hover { background-color: rgb(216, 216, 216); border: 1px solid rgb(198, 198, 198); color: rgb(34, 34, 34); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; }

.ndfHFb-c4YZDc-kODWGd-nK2kYb .ndfHFb-c4YZDc-SxecR { padding-left: 0px !important; padding-right: 2px !important; }

.ndfHFb-c4YZDc-kODWGd-nK2kYb .ndfHFb-c4YZDc-SxecR-skjTt-MFS4be { border-radius: 8px 0px 0px 8px !important; padding-left: 0px !important; padding-right: 3px !important; }

.ndfHFb-c4YZDc-TL3Ynd-V67aGc-haAclf { display: inline-block; }

.ndfHFb-c4YZDc-TL3Ynd-V67aGc { cursor: pointer; display: flex; margin-left: 16px; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-haAclf { display: block; position: absolute; white-space: normal; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b { margin-left: 16px; top: 11px; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-L6cTce { visibility: hidden; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe { border-radius: 24px; height: 24px; padding: 12px; width: 24px; z-index: 101; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe:hover { background: rgb(241, 243, 244); }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe:active { background: rgb(218, 220, 224); }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe { align-items: center; border-radius: 2px; color: rgb(26, 115, 232); display: flex; font-size: 14px; height: 36px; letter-spacing: 0.15px; margin: 6px 0px; min-width: 60px; outline: transparent solid 1px; padding: 0px 15px; z-index: 101; }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe:hover { background: rgb(232, 240, 254); }

.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe:active { background: rgb(210, 227, 252); }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar { height: 12px; overflow: visible; width: 12px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar { width: 16px; }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-button { height: 0px; width: 0px; }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-corner { background: transparent; }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-track { background-color: transparent; border: none; box-shadow: none !important; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track { background-color: rgba(255, 255, 255, 0.1); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track { background: transparent; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-thumb { background-color: rgba(255, 255, 255, 0.9); }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track { background-color: rgba(0, 0, 0, 0.1); }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-thumb { background-color: rgba(0, 0, 0, 0.6); }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb { background-color: rgb(76, 76, 76); background-clip: padding-box; border-style: solid; border-color: transparent; border-width: 0px 1px 0px 0px; box-shadow: rgb(103, 103, 103) 1px 1px 0px inset, rgb(103, 103, 103) 0px -1px 0px inset; min-height: 75px; padding: 100px 0px 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb { background-color: rgba(255, 255, 255, 0.75); border-radius: 1px; border-width: 0px; box-shadow: none; min-height: 56px; padding: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb { background-color: var(--dt-outline-variant,#dadce0); border-radius: 100px; border: 4px solid transparent; background-clip: padding-box; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb { background-color: rgba(0, 0, 0, 0.5); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-to915::-webkit-scrollbar-thumb { background-color: rgb(76, 76, 76); }

.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover { background-color: rgb(159, 159, 159); box-shadow: rgb(204, 204, 204) 1px 1px 0px inset; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover { background-color: rgba(255, 255, 255, 0.9); box-shadow: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover { background-color: var(--dt-outline-variant,#dadce0); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-to915::-webkit-scrollbar-thumb:hover { background-color: rgb(159, 159, 159); }

.ndfHFb-c4YZDc-s2gQvd { }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar { display: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-cYSp0e-s2gQvd.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-track-piece:start { margin-top: 64px; }

.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-uWtm3-ORHb { display: none; align-items: center; background-color: rgb(249, 171, 0); border-radius: 0px; color: rgb(32, 33, 36); height: 3rem; position: relative; top: 0px; width: 100%; z-index: 3; }

.ndfHFb-c4YZDc-uWtm3-ORHb.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb { background: rgb(255, 223, 153); }

.ndfHFb-c4YZDc-uWtm3-ORHb-bN97Pc { align-items: center; display: flex; justify-content: space-between; width: 100%; }

.ndfHFb-c4YZDc-uWtm3-ORHb-Ne3sFf { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-uWtm3-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -1240px; height: 24px; margin: 0px 25px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-Bz112c { margin: 0px 16px; }

.ndfHFb-c4YZDc-uWtm3-ORHb-LQLjdd { display: flex; align-items: center; margin: 8px 0px; order: 0; }

.ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3570px; height: 20px; margin: 0px 25px; width: 20px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-Bz112c { margin: 0px 16px; height: 20px; width: 24px; }

.ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe, .ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe { align-self: center; color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; padding: 0px 8px; text-align: center; text-decoration: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); padding: 0px 12px; }

.ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe:hover, .ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-wvGCSb-gkA7Yd { right: -50px; position: absolute; width: 49px; top: 0px; z-index: 3; }

.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { display: none; }

.ndfHFb-c4YZDc-VCkuzd { min-height: 190px; width: 500px; bottom: 10px; position: absolute; right: 10px; z-index: 10; box-shadow: rgba(0, 0, 0, 0.8) 0px 0px 20px; background-color: rgb(255, 255, 255); padding: 10px; }

.ndfHFb-c4YZDc-VCkuzd::after { content: ""; height: 0px; width: 0px; bottom: -18px; right: 5%; position: absolute; border-top: 18px solid rgb(255, 255, 255); border-left: 15px solid transparent; border-right: 15px solid transparent; }

.ndfHFb-c4YZDc-eLiUMc-Tswv1b-haAclf { margin-bottom: 6px; margin-right: 6px; vertical-align: top; }

.ndfHFb-c4YZDc-eLiUMc-Tswv1b { color: rgb(119, 119, 119); font-size: 8px; }

.ndfHFb-c4YZDc-eLiUMc-Tswv1b-haAclf.ndfHFb-c4YZDc-eLiUMc-Tswv1b { display: flex; position: absolute; right: 0px; bottom: 0px; z-index: 200; }

.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd { border-radius: 2px; border: 0px solid rgb(240, 195, 109); box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; display: none; height: 0px; visibility: hidden; font-size: 11px; overflow: hidden; padding: 0px; text-align: center; background-color: rgb(249, 237, 190); color: rgb(51, 51, 51); }

.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-TSZdd { transition: opacity 0.218s ease 0s; border-width: 1px; display: inline-block; height: auto; max-width: 90%; padding: 6px 16px; text-overflow: ellipsis; visibility: visible; }

.ndfHFb-c4YZDc-X3SwIb.ndfHFb-c4YZDc-b3rLgd-haAclf { height: 0px; position: absolute; text-align: center; top: 50px; width: 100%; z-index: 4; }

.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd { padding-left: 6px; }

.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd, .ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd, .ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited, .ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited { color: rgb(0, 0, 255); cursor: pointer; text-decoration: none; }

.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover, .ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover { text-decoration: underline; }

.ndfHFb-c4YZDc-LgbsSe { cursor: default; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe { cursor: pointer; display: inline-block; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-OWB6Me { cursor: default; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b { background: rgba(66, 133, 244, 0.9); border-color: transparent; border-radius: 50%; border-style: solid; border-width: 30px; display: flex; flex-direction: column; height: 320px; justify-content: center; position: absolute; right: -25px; top: -72px; white-space: normal; width: 320px; z-index: 10; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b-bBybbf { height: 100%; width: 100%; position: relative; z-index: 10; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b .ndfHFb-c4YZDc-jNm5if-Hn6s1b-tJHJj { font-size: 20px; font-weight: normal; line-height: 24px; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b .ndfHFb-c4YZDc-jNm5if-Hn6s1b-Ne3sFf { font-size: 14px; line-height: 24px; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe { position: absolute; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe-Bz112c { background-position: 0px -1632px; height: 24px; left: 32px; opacity: 0.6; position: relative; top: 34px; width: 24px; }

.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe-LkdAo { background: white; border-radius: 50%; height: 88px; left: -32px; position: absolute; top: -34px; width: 88px; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b { animation: 0.6s ease 0s 1 normal none running expandCallout; border-radius: 50%; color: white; justify-content: center; line-height: 24px; position: absolute; transition: all 0s ease-out 0s; white-space: normal; }

@keyframes expandCallout { 
  0% { transform: scale(0, 0); }
  100% { transform: scale(1, 1); }
}

@-webkit-keyframes expandCallout { 
  0% { transform: scale(0, 0); }
  100% { transform: scale(1, 1); }
}

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b-bBybbf { height: 100%; position: relative; width: 100%; z-index: 2; }

.UMrnmb-v3pZbf .ndfHFb-c4YZDc-FNFY6c-Hn6s1b { box-shadow: rgba(17, 109, 231, 0.96) 0px 100px 0px 250px; }

.UMrnmb-nllRtd .ndfHFb-c4YZDc-FNFY6c-Hn6s1b { box-shadow: rgba(21, 138, 54, 0.96) 0px 100px 0px 250px; }

.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-FNFY6c-Hn6s1b { box-shadow: rgba(249, 168, 0, 0.96) 0px 100px 0px 250px; color: black; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-bN97Pc { background-color: rgba(0, 0, 0, 0.004); border: 1px solid transparent; padding: 0px 30px 30px; width: 400px; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-tJHJj { font-size: 20px; font-weight: normal; margin-bottom: 10px; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-Ne3sFf { font-size: 14px; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-KY1xSc-z5C9Gb { color: white; display: inline-block; font-size: 14px; font-weight: bold; margin-left: 10px; text-decoration: none; }

.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-KY1xSc-z5C9Gb { color: black; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-c6xFrd { font-size: 14px; font-weight: bold; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-iDjqhe-Hnhb3b-WtFGnf { border: 1px solid transparent; display: inline-block; }

.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-F2rEXb { border: 1px solid transparent; display: inline-block; margin-left: 40px; opacity: 0.75; }

.UMrnmb-v3pZbf .ndfHFb-c4YZDc-G0brRe-Hn6s1b { background-color: rgba(17, 109, 231, 0.96); }

.UMrnmb-nllRtd .ndfHFb-c4YZDc-G0brRe-Hn6s1b { background-color: rgba(21, 138, 54, 0.96); }

.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b { background-color: rgba(249, 168, 0, 0.96); color: black; }

.ndfHFb-c4YZDc-G0brRe-Hn6s1b { border-radius: 4px 0px 0px 4px; height: 40px; margin: 0px auto; position: absolute; right: 0px; top: 56px; }

.ndfHFb-c4YZDc-G0brRe-Hn6s1b-Ne3sFf { float: left; font-size: 14px; line-height: 40px; margin-bottom: 0px; margin-top: 0px; padding: 0px 32px 0px 24px; }

.ndfHFb-c4YZDc-G0brRe-Hn6s1b-scrj1b-G0brRe { color: white; font-size: 14px; font-weight: bold; line-height: 40px; margin-bottom: 0px; margin-top: 0px; }

.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b-scrj1b-G0brRe { color: black; }

.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b-TvD9Pc { background-position: 0px -1120px; }

.ndfHFb-c4YZDc-G0brRe-Hn6s1b-TvD9Pc { background-position: 0px -3178px; float: right; height: 20px; margin-left: 32px; margin-right: 24px; margin-top: 8px; opacity: 0.5; width: 20px; }

.ndfHFb-c4YZDc-K9a4Re-nKQ6qf { position: absolute; top: 0px; bottom: 0px; width: 100%; user-select: none; }

.ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-oKVyEf { user-select: text; }

.ndfHFb-c4YZDc-MZArnb-b0t70b { box-sizing: border-box; box-shadow: rgb(0, 0, 0) 0px 0px 10px inset; background-color: rgb(36, 34, 35); bottom: 0px; position: fixed; right: 0px; top: 47px; width: 400px; z-index: 1; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b { box-shadow: none; background-color: rgb(50, 50, 50); width: 344px; top: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b { background: none; padding: 0px 16px 16px 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b-haAclf { background: var(--dt-surface,#fff); border-radius: 24px; height: 100%; display: flex; flex-direction: column; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b { z-index: 4; }

.ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce { display: none; }

.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c { display: block; margin-left: auto; margin-right: auto; }

.ndfHFb-c4YZDc-MZArnb-tJHJj { box-sizing: border-box; font-family: Roboto, arial, sans-serif; font-size: 14px; text-transform: uppercase; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj { box-shadow: rgba(0, 0, 0, 0.3) 0px 2px 2px; font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 16px; text-transform: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj { box-shadow: none; border-bottom: solid 2px var(--dt-outline-variant,#dadce0); }

.ndfHFb-c4YZDc-MZArnb-bN97Pc { inset: 50px 0px 0px; margin: 5px 0px; overflow-y: auto; position: absolute; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MZArnb-bN97Pc { position: static; top: 0px; margin: 5px 0px 15px; }

.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e { box-sizing: border-box; color: rgb(192, 190, 190); cursor: pointer; display: inline-block; height: 50px; line-height: 50px; margin: 0px 16px; padding: 4px 2px 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e { height: 56px; line-height: 56px; }

.ndfHFb-c4YZDc-MZArnb-cXCLoc { border-bottom: 1px solid rgb(204, 204, 204); margin: 0px 15px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-cXCLoc { border-bottom: none; display: inline-block; margin: 0px; }

.ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd.ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge { border-bottom: 3px solid rgb(77, 144, 254); }

.ndfHFb-c4YZDc-MZArnb-AznF2e:hover.ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge { border-bottom: 3px solid rgb(100, 100, 100); }

.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e:hover { margin: 0px 18px; padding: 4px 0px 0px; }

.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e.ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd { color: rgb(255, 255, 255); cursor: default; }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj { color: rgb(238, 238, 238); font-family: Roboto-light, arial, sans-serif; height: 40px; line-height: 40px; }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS { background-color: rgb(36, 34, 35); float: left; font-family: Roboto-light, arial, sans-serif; font-size: 12px; font-weight: 500; padding-right: 5px; text-transform: uppercase; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS { background-color: rgb(50, 50, 50); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; text-transform: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS { background: var(--dt-surface,#fff); }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf { margin-bottom: 10px; padding-top: 19px; width: 100%; }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe { border-top: 1px solid rgb(104, 104, 104); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe { border-top: 1px solid rgba(255, 255, 255, 0.15); }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc { color: rgb(182, 182, 182); font-size: 12px; padding-bottom: 20px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc { color: rgba(255, 255, 255, 0.57); }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b { display: inline-block; text-align: left; width: calc(100% - 150px); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b { color: rgba(255, 255, 255, 0.9); width: calc(100% - 128px); }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc { display: inline-block; }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc { vertical-align: top; width: 150px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc { width: 128px; }

.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-BA389-V67aGc { width: calc(100% - 100px); }

.ndfHFb-c4YZDc-MZArnb-P86uke-PntVL { display: inline-block; vertical-align: top; width: 100%; }

.ndfHFb-c4YZDc-MZArnb-P86uke-Bz112c { float: left; margin-right: 12px; margin-top: 5px; width: 16px; height: 13px; }

.ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd { cursor: pointer; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd:focus, .ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd:hover { text-decoration: underline; }

.ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d { line-height: 24px; margin-left: 36px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.ndfHFb-c4YZDc-MZArnb-BA389-nNAX0 { display: inline-block; float: right; overflow-x: hidden; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BA389-nNAX0 { color: rgba(255, 255, 255, 0.9); }

.ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c { line-height: 24px; padding-bottom: 10px; }

.ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc { box-sizing: content-box; border: none; width: 100%; }

.ndfHFb-c4YZDc-MZArnb-ij8cu { font-weight: normal; padding-bottom: 20px; overflow-wrap: break-word; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-ij8cu { margin-right: 44px; }

.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe { background-color: rgb(36, 34, 35); cursor: pointer; float: right; margin-top: 8px; padding-left: 3px; }

.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgb(36, 34, 35); background-image: -webkit-linear-gradient(top, rgb(51, 51, 51), rgb(34, 34, 34)); }

.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -760px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-MZArnb-ij8cu-DyVDA { box-sizing: border-box; min-height: 75px; max-width: 350px; overflow-y: auto; width: 100%; }

.ndfHFb-c4YZDc-MZArnb-Tswv1b-nUpftc, .ndfHFb-c4YZDc-MZArnb-RDNXzf-nUpftc { user-select: text; padding: 15px; }

.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS { font-size: 12px; line-height: 20px; }

.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c { margin: 1px 0px; }

.ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c { float: left; height: 24px; }

.ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c .ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c { height: 24px; position: relative; width: 24px; }

.ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e { background-color: rgb(70, 68, 69); border-radius: 50%; display: inline-block; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb { color: rgb(255, 255, 255); line-height: 24px; text-align: center; text-transform: uppercase; vertical-align: middle; }

.ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c { background-position: 0px -2160px; }

.ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c { background-position: 0px -2400px; }

.ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c-SfQLQb-hSRGPd { background-position: 0px -280px; }

.ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c { background-position: 0px -720px; }

.ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c-SfQLQb-hSRGPd { background-position: 0px -480px; }

.ndfHFb-c4YZDc-MZArnb-YLEF4c-Bz112c { height: 20px; margin: 2px; width: 20px; }

.ndfHFb-c4YZDc-MZArnb-nupQLb-BA389-Ne3sFf { display: inline-block; }

.ndfHFb-c4YZDc-MZArnb-MPu53c { box-sizing: border-box; border: 2px solid rgb(193, 191, 191); border-radius: 2px; cursor: pointer; float: right; height: 20px; width: 20px; }

.ndfHFb-c4YZDc-MZArnb-MPu53c-bN97Pc { height: 16px; }

.ndfHFb-c4YZDc-MZArnb-MPu53c-fmcmS { font-size: 20px; font-weight: bold; line-height: 16px; position: absolute; }

.ndfHFb-c4YZDc-MZArnb-MPu53c-Bz112c { background-position: 0px -1680px; display: inline-block; height: 14px; width: 14px; margin-top: 2px; margin-left: 1px; }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b { width: 100%; right: 0px; transition: right 0.218s cubic-bezier(0, 0, 0.2, 1) 0s; }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce { display: block; right: -100%; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -288px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-J2xVie-Bz112c { background-position: 0px -3674px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c { background-position: 0px -3138px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c { background-position: 0px -1264px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c-SfQLQb-hSRGPd { background-position: 0px -816px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c { background-position: 0px -168px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c-SfQLQb-hSRGPd { background-position: 0px -736px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe:not(.ndfHFb-c4YZDc-LgbsSe-ZmdkE) { background-color: rgb(50, 50, 50); padding: 8px; margin-top: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe:not(.ndfHFb-c4YZDc-LgbsSe-ZmdkE) { background-color: transparent; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe { background-color: rgba(196, 199, 197, 0.12); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { float: right; margin: 8px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -3178px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { margin-top: -8px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb { border-top: 1px solid rgb(104, 104, 104); font-size: 12px; font-weight: normal; outline: none; padding: 18px 0px 7px; position: relative; zoom: 1; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb:first-child { border-top-color: transparent; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-haAclf { margin-left: 55px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if { min-height: 48px; position: relative; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-tJHJj { color: rgb(117, 114, 114); font-style: italic; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-EieU8 { background-color: rgb(33, 31, 32); margin: 4px 0px 3px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb { margin-bottom: 10px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od { color: rgb(182, 182, 182); display: inline-block; font-weight: bold; max-width: 180px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-IIEkAe .ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od { max-width: 120px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc .ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od { font-style: normal; margin-right: 4px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c { border-radius: 50%; height: 48px; left: 0px; position: absolute; width: 48px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c { border-radius: 0px; height: 24px; left: 6px; width: 24px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e { height: 48px; width: 48px; left: 0px; position: absolute; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb { font-size: 24px; line-height: 48px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e { border-radius: 0px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb { font-size: 12px; line-height: 24px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb-haAclf { color: rgb(193, 191, 191); font-size: 10px; padding-top: 2px; position: absolute; right: 0px; top: 0px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb { display: inline-block; padding: 0px 3px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc .ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb { color: rgb(193, 191, 191); font-size: 10px; padding: 3px 0px; position: relative; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-bN97Pc { color: rgb(255, 255, 255); margin-top: 5px; overflow-wrap: break-word; top: -7px; zoom: 1; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb { border-top: 1px solid rgb(36, 34, 35); color: rgb(136, 136, 136); min-height: 24px; padding: 6px 3px 0px 6px; position: relative; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb:first-child { border-top-color: transparent; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc { padding-left: 30px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-fmcmS { line-height: 140%; position: relative; top: -3px; width: 100%; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-qJTHM { color: rgb(255, 255, 255); display: inline; margin: 0px; position: relative; top: -4px; width: 100%; overflow-wrap: break-word; }

.ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Ne3sFf { display: inline; padding-right: 18px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-JIbuQc { color: rgb(255, 255, 255); display: inline; font-style: italic; position: relative; top: -4px; }

.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-JIbuQc + .ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-qJTHM { display: block; }

.ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Bz112c { background-position: 0px -1680px; display: inline-block; height: 12px; margin-left: 3px; position: absolute; right: 0px; width: 15px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Bz112c { background-position: 0px -2504px; }

.ndfHFb-c4YZDc-C7uZwb-LgbsSe .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { opacity: 0.87; margin-left: auto; margin-right: auto; margin-top: 3px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { opacity: 0.87; margin-right: auto; margin-top: 3px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c.ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { opacity: 0.47; }

.ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-nupQLb-Bz112c { background-position: 0px -1040px; }

.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c { background-position: 0px -1880px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c { background-position: 0px -1560px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c { background-position: 0px -2480px; }

.ndfHFb-c4YZDc-VkLyEc-Bz112c { background-position: 0px -2320px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c { background-position: 0px -1480px; }

.ndfHFb-c4YZDc-euCgFf-Bz112c { background-position: 0px -1440px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c { background-position: 0px -1200px; }

.ndfHFb-c4YZDc-hN7jy-Bz112c { background-position: 0px -2200px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c { background-position: 0px -2280px; }

.ndfHFb-c4YZDc-PEFSMe-Bz112c { background-position: 0px -2240px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c { background-position: 0px -360px; }

.ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c { background-position: 0px -1800px; }

.ndfHFb-c4YZDc-w37qKe-Bz112c { background-position: 0px -440px; }

.ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c { background-position: 0px -40px; }

.ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c { background-position: 0px -1720px; }

.ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c { background-position: 0px -2000px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg"); background-size: auto; margin-left: 2px; left: 8px; top: 3px; }

.ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { top: 2px; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c.ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c, .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c.ndfHFb-c4YZDc-w37qKe-Bz112c { height: 24px; margin-left: 0px; margin-top: -1px; width: 24px; }

.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe { border: 1px solid rgb(26, 115, 232); border-radius: 2px; box-shadow: rgba(101, 101, 101, 0.1) 0px 1px 0px inset; background-color: rgb(26, 115, 232); color: rgb(255, 255, 255); display: inline-block; font-size: 11px; font-weight: bold; text-align: center; text-shadow: rgba(0, 0, 0, 0.8) 0px 1px 0px; height: 28px; line-height: 28px; margin-top: 20px; min-width: 54px; padding: 0px 20px 0px 7px; vertical-align: middle; white-space: nowrap; }

.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg"); height: 21px; margin-top: 4px; position: absolute; width: 21px; }

.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-fmcmS { margin-left: 35px; margin-right: 10px; }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe { background-color: rgb(26, 115, 232); background-image: -webkit-linear-gradient(top, rgb(26, 115, 232), rgb(53, 122, 232)); }

.ndfHFb-c4YZDc-LgbsSe-auswjd.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe { box-shadow: rgba(0, 0, 0, 0.8) 0px 1px 6px inset; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-C7uZwb-LgbsSe .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { margin-top: 0px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { margin-top: 0px; height: 24px; width: 24px; background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nupQLb-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nupQLb-Bz112c { background-position: 0px -2384px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c { background-position: 0px -408px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c { background-position: 0px -3530px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c { background-position: 0px -408px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c { background-position: 0px -2384px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c { background-position: 0px -632px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-VkLyEc-Bz112c { background-position: 0px -2584px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c { background-position: 0px -2890px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-VkLyEc-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c { background-position: 0px -2584px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-euCgFf-Bz112c { background-position: 0px -3218px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c { background-position: 0px -2994px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-euCgFf-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c { background-position: 0px -3218px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hN7jy-Bz112c { background-position: 0px -2016px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c { background-position: 0px -1368px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hN7jy-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c { background-position: 0px -2016px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c { background-position: 0px -3258px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c { background-position: 0px -1856px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c { background-position: 0px -3258px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-PEFSMe-Bz112c { background-position: 0px -3426px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c { background-position: 0px -512px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-PEFSMe-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c { background-position: 0px -3426px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c { background-position: 0px -3098px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c { background-position: 0px -3714px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-w37qKe-Bz112c { background-position: 0px -1200px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-w37qKe-Bz112c { background-position: 0px -1568px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c { background-position: 0px -672px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c { background-position: 0px -328px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c { background-position: 0px -2930px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c { background-position: 0px -1672px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c { background-position: 0px -88px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c { background-position: 0px -1488px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-Bz112c { background-position: 0px -1712px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-Bz112c { background-position: 0px -208px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-GSQQnc-LgbsSe { background-position: 0px -368px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-GSQQnc-LgbsSe { background-position: 0px -2304px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c { background-position: 0px -2602px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3338px; transform: scale(0.8) translateX(3px) translateY(9px); width: 24px; height: 24px; pointer-events: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-hOcTPc .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c { transform: scale(0.8); margin-left: 4px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-RDNXzf-OWB6Me-Bz112c { background-position: 0px -40px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c { background-position: 0px -1632px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c { background-position: 0px -2602px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ge6pde-Bz112c .ndfHFb-aZ2wEe { display: block; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-pGuBYc-Bz112c { background-position: 0px -472px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-MqcBrc-Bz112c { background-position: 0px -3634px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-MqcBrc-Bz112c { background-position: 0px -2850px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-SjW3R-Bz112c { background-position: 0px -3034px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-SjW3R-Bz112c { background-position: 0px -2970px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-lCdvJf-Bz112c { background-position: 0px -1896px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-lCdvJf-Bz112c { background-position: 0px -128px; }

.ndfHFb-c4YZDc-E90Ek { background-color: rgba(0, 0, 0, 0.75); display: inline-block; margin-right: 50px; padding: 2px; width: 500px; }

.ndfHFb-c4YZDc-E90Ek-tJHJj { font-size: 18px; margin: 10px; text-align: center; }

.ndfHFb-c4YZDc-E90Ek-LgbsSe { background-color: dimgray; cursor: pointer; float: right; padding: 10px; }

.ndfHFb-c4YZDc-E90Ek-bN97Pc { max-height: 600px; max-width: 600px; overflow-x: scroll; }

.ndfHFb-c4YZDc-E90Ek-Tswv1b-tJHJj { margin: 10px; text-align: left; }

.ndfHFb-c4YZDc-E90Ek-Tswv1b-lTBxed { color: white; margin: 0px 10px; }

.ndfHFb-c4YZDc-Sx9Kwc { background: padding-box rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.333); box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; outline: 0px; padding: 30px 42px; position: absolute; z-index: 102; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-Sx9Kwc { background: var(--dt-surface,#fff); padding: 24px; border-radius: 8px; }

.ndfHFb-c4YZDc-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); left: 0px; position: absolute; top: 0px; z-index: 101; }

.ndfHFb-c4YZDc-qbOKL-OEVmcd .VIpgJd-TUo6Hb-xJ5Hnf, .ndfHFb-c4YZDc-qbOKL-OEVmcd .XKSfm-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); }

div.ndfHFb-c4YZDc-Sx9Kwc-xJ5Hnf { opacity: 0.75; }

.ndfHFb-c4YZDc-Sx9Kwc-r4nke { background-color: rgb(255, 255, 255); color: rgb(0, 0, 0); cursor: default; font-size: 16px; line-height: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-r4nke { background-color: var(--dt-surface,#fff); color: var(--dt-on-surface,#3c4043); font: var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-headline-small-spacing,0); }

.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc { height: 11px; opacity: 0.7; padding: 17px; position: absolute; right: 0px; top: 0px; width: 11px; }

.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc::after { content: ""; background: url("//ssl.gstatic.com/ui/v1/dialog/close-x.png"); position: absolute; height: 11px; width: 11px; right: 17px; }

.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.ndfHFb-c4YZDc-Sx9Kwc-bN97Pc { background-color: rgb(255, 255, 255); line-height: 1.4em; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-bN97Pc { background-color: var(--dt-surface,#fff); }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button { border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); cursor: default; font-size: 11px; font-weight: bold; height: 29px; line-height: 27px; margin: 0px 16px 0px 0px; min-width: 72px; outline: 0px; padding: 0px 8px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button { margin: 0px 0px 0px 24px; border-radius: 100px; background: var(--dt-surface,#fff); color: var(--dt-primary,#1a73e8); font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); border: none; }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:hover, .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:hover { background: rgba(168, 199, 250, 0.08); color: var(--dt-primary,#1a73e8); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active { background: rgba(168, 199, 250, 0.12); color: var(--dt-primary,#1a73e8); border: none; outline: none; box-shadow: none; }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:focus { border: 1px solid rgb(77, 144, 254); }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button[disabled] { box-shadow: none; background: none rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc { background-color: rgb(26, 115, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(71, 135, 237)); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:hover { background-color: rgb(53, 122, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:active { background-color: rgb(53, 122, 232); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc[disabled] { box-shadow: none; background: rgb(77, 144, 254); color: rgb(255, 255, 255); opacity: 0.5; }

.ndfHFb-c4YZDc-Sx9Kwc-TD02Lb { position: absolute; visibility: hidden; }

.ndfHFb-c4YZDc-uoC0bf .XKSfm-Sx9Kwc { padding: 24px; border-radius: 0.5rem; }

.ndfHFb-c4YZDc-uoC0bf .XKSfm-Sx9Kwc-r4nke { font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 24px; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe { display: flex; align-items: center; position: absolute; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-B8qYne, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-B8qYne, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-B8qYne { height: 100%; width: 100%; display: none; align-items: center; position: absolute; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-B8qYne-RJLb9c, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-B8qYne-RJLb9c, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-B8qYne-RJLb9c { max-width: 100%; max-height: 100%; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-WbpZL, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-WbpZL, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-WbpZL { height: 100%; width: 100%; display: none; align-items: center; z-index: 2; pointer-events: all; background: rgb(232, 240, 254); color: rgb(24, 90, 188); border: 1px solid rgb(24, 90, 188); border-radius: 4px; box-sizing: border-box; cursor: pointer; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-jf2N7b-dIxMhd-zUk4Qd, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-jf2N7b-dIxMhd-zUk4Qd, .ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-jf2N7b-dIxMhd-zUk4Qd, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-jf2N7b-dIxMhd-zUk4Qd { height: 100%; width: 100%; display: none; align-items: center; z-index: 2; pointer-events: all; background: rgb(241, 243, 244); color: rgb(192, 192, 192); border: 1px solid rgb(192, 192, 192); border-radius: 4px; box-sizing: border-box; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-jf2N7b-dIxMhd-MFS4be, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-jf2N7b-dIxMhd-MFS4be, .ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-jf2N7b-dIxMhd-MFS4be, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-jf2N7b-dIxMhd-MFS4be { height: 100%; width: 100%; display: none; align-items: center; z-index: 2; pointer-events: all; background: transparent; color: rgb(192, 192, 192); border: 1px solid rgb(192, 192, 192); border-radius: 4px; box-sizing: border-box; }

.ndfHFb-c4YZDc-dZssN-yrriRe-JbbQac-LgbsSe { position: absolute; right: 0px; top: 0px; background: rgb(60, 64, 67); opacity: 0.4; border-radius: 50%; display: none; height: 24px; width: 24px; pointer-events: all; z-index: 2; cursor: pointer; }

.ndfHFb-c4YZDc-dZssN-yrriRe-JbbQac-LgbsSe-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3362px; height: 11.62px; width: 11.67px; margin: auto; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-WbpZL-fmcmS, .ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-WbpZL-fmcmS, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-WbpZL-fmcmS { color: rgb(23, 78, 166); font-family: "Roboto Mono", monospace; font-style: normal; font-weight: bold; font-size: 16px; line-height: 22px; position: absolute; inset: auto 78% auto 9.41%; }

.ndfHFb-c4YZDc-dZssN-mKZypf-qFWjAd-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -2786px; height: 13.33px; width: 13.29px; position: absolute; top: auto; bottom: auto; right: 14.31%; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe { display: flex; justify-content: center; align-items: center; position: absolute; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-fmcmS { display: none; font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 22px; line-height: 20px; color: black; text-size-adjust: auto; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-suEOdc { position: absolute; background-color: rgb(32, 33, 36); color: rgb(218, 220, 224); font-family: Roboto; font-style: normal; font-weight: 400; font-size: 14px; line-height: 20px; letter-spacing: 0.2px; border-radius: 4px; visibility: hidden; width: 210px; height: max-content; top: 42px; left: 20px; padding: 9px 13px; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe:hover .ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-suEOdc { position: absolute; visibility: visible; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe:hover { z-index: 100; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-FVVVue-WAutxc-zUk4Qd { display: none; width: 100%; height: 100%; align-items: center; background-color: rgb(232, 240, 254); color: rgb(23, 78, 166); position: absolute; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -2136px; height: 17.61px; width: 16px; position: absolute; top: auto; bottom: auto; left: 18.5px; transform: scale(0.9375, 0.9432); }

.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-FVVVue-WAutxc-zUk4Qd, .ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-FVVVue-WAutxc-zUk4Qd, .ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-FVVVue-WAutxc-zUk4Qd { display: none; width: 100%; height: 100%; align-items: center; background-color: rgb(232, 240, 254); color: rgb(23, 78, 166); position: absolute; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -1608px; height: 17.61px; width: 16px; position: absolute; top: auto; bottom: auto; left: 18.5px; transform: scale(0.9375, 0.9432); }

.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3506px; height: 24px; width: 24px; position: absolute; top: auto; bottom: auto; left: 18.5px; transform: scale(0.9375, 0.9432); }

.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -1792px; height: 24px; width: 24px; position: absolute; top: auto; bottom: auto; left: 18.5px; transform: scale(0.9375, 0.9432); }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 453px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc { background: rgb(31, 31, 31); display: inline; width: 444px; }

.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 340px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc { background: rgb(31, 31, 31); display: inline; width: 444px; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 468px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc { background: rgb(31, 31, 31); width: 468px; }

.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 300px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc { background: rgb(31, 31, 31); border-radius: 8px; display: inline; width: 444px; }

.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 350px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc { background: rgb(31, 31, 31); border-radius: 8px; display: inline; width: 444px; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-xJ5Hnf, .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-xJ5Hnf, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-xJ5Hnf, .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-xJ5Hnf, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); height: 100%; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 101; }

.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-xJ5Hnf { background-color: rgb(0, 0, 0); height: 100%; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 101; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke { margin: 0px auto; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke { margin: 24px 24px 0px; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-r4nke, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-r4nke, .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-r4nke, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-r4nke { margin: 24px; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1.375rem; font-weight: 400; letter-spacing: 0px; line-height: 1.75rem; color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-r4nke-fmcmS { color: rgb(197, 199, 197); }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-HiaYvf { width: 125px; height: 125px; margin: 39px auto 33px; display: block; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-HiaYvf { display: none; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-bN97Pc { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; color: rgb(95, 99, 104); display: flex; flex-direction: column; justify-content: space-between; margin: 16px 24px 12px; text-align: center; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-bN97Pc { margin: 12px; color: rgb(197, 199, 197); text-align: left; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-bN97Pc { color: rgb(95, 99, 104); display: flex; flex-direction: column; justify-content: space-between; margin: 0px 12px 12px; text-align: left; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-g7W7Ed { color: rgb(95, 99, 104); font-family: Roboto; font-style: normal; font-weight: 400; font-size: 14px; line-height: 20px; letter-spacing: 0.2px; margin-bottom: 22.6px; width: 428px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-g7W7Ed { color: rgb(197, 199, 197); }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-MPu53c-bN97Pc { color: rgb(60, 64, 67); font-family: Roboto; font-style: normal; font-weight: 700; font-size: 14px; line-height: 20px; letter-spacing: 0.2px; text-align: left; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-MPu53c-bN97Pc { color: rgb(197, 199, 197); font-weight: 400; }

.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-bN97Pc { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; color: rgb(95, 99, 104); display: flex; flex-direction: column; justify-content: space-between; margin: 16px 24px 12px; text-align: center; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-bN97Pc { color: rgb(197, 199, 197); align-items: flex-start; margin: 0px 12px; text-align: left; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-bN97Pc-PLDbbf { text-decoration: none; color: rgb(26, 115, 232); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-bN97Pc-PLDbbf { text-decoration: none; color: rgb(168, 199, 250); }

.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-bN97Pc { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; color: rgb(95, 99, 104); justify-content: space-between; margin: 0px 24px; max-width: 300px; overflow-wrap: break-word; text-align: center; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-bN97Pc { margin: 12px; color: rgb(197, 199, 197); text-align: left; }

.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-bN97Pc { color: rgb(95, 99, 104); display: flex; flex-direction: column; justify-content: space-between; text-align: center; margin: 0px 12px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-bN97Pc { color: rgb(197, 199, 197); align-items: flex-start; margin: 0px 12px; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-LgbsSe, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-LgbsSe, .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-IbE0S-LgbsSe, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-IbE0S-LgbsSe, .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 20px; background: rgb(255, 255, 255); border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(26, 115, 232); margin: 0px 12px; min-width: 70px; outline: none; padding: 8px 24px; text-align: center; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-IbE0S-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-IbE0S-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-LgbsSe { background: transparent; color: rgb(168, 199, 250); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-LgbsSe { background: rgb(168, 199, 250); color: var(--dt-on-primary,#fff); border: none; border-radius: 100px; margin: 0px 18px; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 20px; border: none; background: rgb(26, 115, 232); box-sizing: border-box; border-radius: 4px; color: rgb(255, 255, 255); margin: 0px 12px; min-width: 70px; outline: none; padding: 8px 24px; text-align: center; cursor: pointer; opacity: 0.3; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe { border-radius: 100px; background: rgb(168, 199, 250); color: var(--dt-on-primary,#fff); }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-qnnXGd { opacity: 1; }

.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-ERydpb-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 20px; border: none; background: rgb(217, 48, 37); box-sizing: border-box; border-radius: 4px; color: rgb(255, 255, 255); margin: 0px 12px; min-width: 70px; outline: none; padding: 8px 24px; text-align: center; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-ERydpb-LgbsSe { background: var(--dt-error,#d93025); color: var(--dt-on-primary,#fff); border-radius: 100px; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-HiaYvf { width: 97px; height: 97px; margin-bottom: 36px; margin-right: auto; margin-left: auto; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-HiaYvf { display: none; }

.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-c6xFrd { margin: 21px; display: flex; flex-direction: row; padding: 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-c6xFrd, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-c6xFrd, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-c6xFrd { justify-content: flex-end; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-c6xFrd, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-c6xFrd { margin-left: auto; margin-right: auto; margin-bottom: 18px; display: flex; flex-direction: row; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-c6xFrd { margin-top: 18px; justify-content: flex-end; }

.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-c6xFrd { margin-right: 22px; margin-left: auto; margin-bottom: 18px; display: flex; flex-direction: row; padding: 0px; }

.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-c6xFrd { margin: 22px 22px 18px auto; display: flex; flex-direction: row; padding: 0px; }

.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-IbE0S-LgbsSe .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-ERydpb-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-IbE0S-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-dZssN-ORHb-haAclf { display: none; position: relative; top: 0px; z-index: 3; }

.ndfHFb-c4YZDc-dZssN-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: block; }

.ndfHFb-c4YZDc-dZssN-ORHb { align-items: center; display: flex; letter-spacing: 0.00625em; font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1rem; font-weight: 500; line-height: 1.5rem; background-color: rgb(232, 240, 254); border-radius: 0px; color: rgb(32, 33, 36); height: 48px; width: 100%; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb { background: rgb(168, 199, 250); }

.ndfHFb-c4YZDc-dZssN-ORHb-bN97Pc { align-items: center; display: flex; justify-content: space-between; width: 100%; }

.ndfHFb-c4YZDc-dZssN-ORHb-jOfkMb { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-jOfkMb { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); }

.ndfHFb-c4YZDc-dZssN-ORHb-Vkfede-Ne3sFf { margin-left: 16px; margin-right: auto; font-size: 14px; font-weight: 400; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-Vkfede-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-dZssN-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -712px; height: 16px; margin: 0px 13px 0px 25px; width: 18px; transform: scale(1.076, 1); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-Bz112c { background-position: 0px -976px; height: 24px; margin: 0px 16px; width: 24px; }

.ndfHFb-c4YZDc-dZssN-ORHb-LQLjdd { display: flex; flex: 0 0 auto; -webkit-box-flex: 0; margin: 8px 0px; order: 0; }

.ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe, .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe { color: rgb(26, 115, 232); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; border-radius: 5px; letter-spacing: 0.25px; line-height: 20px; text-align: center; text-decoration: none; margin: 0px 12px; padding: 6px 14px; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe { color: rgb(32, 33, 36); background: transparent; font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); }

.ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe:hover { background: rgb(248, 251, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe:hover { background: transparent; }

.ndfHFb-c4YZDc-dZssN-ORHb-LgbsSe-L6cTce { display: none; }

.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe { color: rgb(255, 255, 255); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; border-radius: 5px; letter-spacing: 0.25px; line-height: 20px; text-align: center; text-decoration: none; margin: 0px 12px; padding: 6px 14px; background-color: rgb(26, 115, 232); cursor: pointer; opacity: 0.3; pointer-events: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe { color: rgb(255, 255, 255); background: var(--dt-on-primary,#fff); font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); opacity: 0.38; border-radius: 100px; }

.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe:hover { background: rgb(43, 125, 233); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe:hover { background: var(--dt-on-primary,#fff); }

.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-sM5MNb, .ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-sM5MNb, .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-sM5MNb { background: none; }

.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe.ndfHFb-c4YZDc-LgbsSe-qnnXGd { opacity: 1; pointer-events: auto; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf { display: none; align-items: center; letter-spacing: 0.00625em; font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1rem; font-weight: 500; line-height: 1.5rem; background-color: rgb(232, 240, 254); border-radius: 0px; color: rgb(32, 33, 36); height: 48px; width: 100%; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf { background: rgb(168, 199, 250); }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-bN97Pc { align-items: center; display: flex; justify-content: space-between; width: 100%; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-jOfkMb { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-jOfkMb { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Vkfede-Ne3sFf { margin-left: 16px; margin-right: auto; font-size: 14px; font-weight: 400; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Vkfede-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -712px; height: 16px; margin: 0px 13px 0px 25px; width: 18px; transform: scale(1.076, 1); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Bz112c { background-position: 0px -976px; height: 24px; margin: 0px 16px; width: 24px; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-LQLjdd { display: flex; flex: 0 0 auto; -webkit-box-flex: 0; margin: 8px 0px; order: 0; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe, .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe { color: rgb(26, 115, 232); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; border-radius: 5px; letter-spacing: 0.25px; line-height: 20px; text-align: center; text-decoration: none; margin: 0px 12px; padding: 6px 14px; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-mKZypf-LgbsSe { color: rgb(32, 33, 36); background: transparent; font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe:hover, .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe:hover { background: rgb(248, 251, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-mKZypf-LgbsSe:hover { background: transparent; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe { color: rgb(255, 255, 255); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; border-radius: 5px; letter-spacing: 0.25px; line-height: 20px; text-align: center; text-decoration: none; margin: 0px 12px; padding: 6px 14px; background-color: rgb(26, 115, 232); cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe { border-radius: 100px; background: var(--dt-on-primary,#fff); cursor: pointer; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe:hover { background: rgb(43, 125, 233); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe:hover { background: var(--dt-on-primary,#fff); }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-sM5MNb, .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-sM5MNb, .ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-sM5MNb { background: none; }

.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-dZssN-x5yx9d-b0t70b { background: white; bottom: 0px; position: absolute; right: 0px; top: 0px; display: none; }

.ndfHFb-c4YZDc-dZssN-x5yx9d-L5Fo6c { border: none; height: 100%; width: 100%; }

.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe { width: 100%; height: 100%; top: 50%; }

.ndfHFb-c4YZDc-EglORb-ge6pde.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe { min-width: 0px; }

.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-haAclf { z-index: 9000; }

.ndfHFb-c4YZDc-dZssN-G0KQoc { position: absolute; width: 100%; height: 100%; z-index: 2; pointer-events: all; }

.ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c { background-repeat: no-repeat; opacity: 0.87; margin-left: auto; margin-right: auto; margin-top: 3px; height: 21px; width: 19px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-PlOyMe-bN97Pc { line-height: 32px; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-spinner_dark.gif"); }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-Wrql6b-PlOyMe { background-color: transparent; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: none; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: none; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c .ndfHFb-aZ2wEe { display: block; }

.ndfHFb-c4YZDc-cnqxLd { background-color: rgb(18, 18, 18); bottom: 0px; color: rgb(255, 255, 255); font-size: 0px; height: 0px; position: absolute; transition: height 0.218s ease-out 0s; width: 100%; z-index: 2; }

.ndfHFb-c4YZDc-cnqxLd-SmKAyb { overflow: auto hidden; position: absolute; top: 0px; width: 100%; white-space: nowrap; }

.ndfHFb-c4YZDc-cnqxLd-OEVmcd { border: 3px solid rgb(255, 255, 255); border-radius: 3px; position: absolute; height: 63px; width: 84px; margin-top: 3px; }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd { position: absolute; height: 25px; z-index: 1; }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd-hOcTPc { left: 12px; }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd-AeOLfc { right: 12px; }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe { background-color: rgba(0, 0, 0, 0.2); border-radius: 3px; color: rgba(255, 255, 255, 0.87); font-size: 11px; text-align: center; text-shadow: rgba(0, 0, 0, 0.8) 0px 1px 1px; height: 25px; line-height: 25px; padding: 0px 13px; }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgba(0, 0, 0, 0.4); }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-IwzHHe, .ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-cnqxLd-N7Eqid-bF1uUb { background-color: rgba(0, 0, 0, 0.6); }

.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE, .ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-cnqxLd-N7Eqid-bF1uUb.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgba(0, 0, 0, 0.9); }

.ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c { background-position: 0px -1080px; display: inline-block; height: 21px; margin-right: 4px; vertical-align: top; width: 21px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c { background-position: 0px -2160px; }

.ndfHFb-c4YZDc-cnqxLd-LSZ0mb.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c { background-position: 0px -960px; height: 16px; margin-top: 5px; padding-left: 5px; width: 16px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cnqxLd-LSZ0mb.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c { background-position: 0px -1936px; }

.ndfHFb-c4YZDc-cnqxLd-LSZ0mb-fmcmS { display: inline-block; margin-top: 1px; vertical-align: middle; }

.ndfHFb-c4YZDc-n5VRYe-ma6Yeb, .ndfHFb-c4YZDc-n5VRYe-AeOLfc, .ndfHFb-c4YZDc-n5VRYe-cGMI2b, .ndfHFb-c4YZDc-n5VRYe-hOcTPc { z-index: 1; position: absolute; }

.ndfHFb-c4YZDc-n5VRYe-ma6Yeb, .ndfHFb-c4YZDc-n5VRYe-cGMI2b { height: 8px; left: 0px; right: 0px; }

.ndfHFb-c4YZDc-n5VRYe-AeOLfc, .ndfHFb-c4YZDc-n5VRYe-hOcTPc { bottom: 0px; top: 0px; width: 8px; }

.ndfHFb-c4YZDc-n5VRYe-ma6Yeb { background-image: -webkit-linear-gradient(top, rgba(0, 0, 0, 0.35), rgba(0, 0, 0, 0)); top: 0px; }

.ndfHFb-c4YZDc-n5VRYe-AeOLfc { background-image: -webkit-linear-gradient(right, rgba(0, 0, 0, 0.35), rgba(0, 0, 0, 0)); right: 0px; }

.ndfHFb-c4YZDc-n5VRYe-cGMI2b { background-image: -webkit-linear-gradient(bottom, rgba(0, 0, 0, 0.35), rgba(0, 0, 0, 0)); bottom: 0px; }

.ndfHFb-c4YZDc-n5VRYe-hOcTPc { background-image: -webkit-linear-gradient(left, rgba(0, 0, 0, 0.35), rgba(0, 0, 0, 0)); left: 0px; }

.ndfHFb-c4YZDc-Sx9Kwc.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc { padding: 0px; }

.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde { background-color: rgb(243, 243, 243); height: 100%; position: relative; width: 100%; }

.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde .ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde-k4Qmrd { text-align: center; width: 100%; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-ge6pde-RJLb9c { background-image: url("//ssl.gstatic.com/ui/v1/activityindicator/loading_bg_f5.gif"); background-repeat: no-repeat; display: inline-block; height: 19px; position: relative; top: 3px; width: 19px; }

.ndfHFb-c4YZDc-w5vlXd { border: 1px solid transparent; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited) { background-repeat: no-repeat; background-image: url("//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg") !important; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg") !important; }

.ndfHFb-c4YZDc-L5Fo6c-nUpftc { position: absolute; }

.ndfHFb-c4YZDc-HiaYvf { position: absolute; background-color: white; background-image: linear-gradient(45deg, rgb(239, 239, 239) 25%, transparent 25%, transparent 75%, rgb(239, 239, 239) 75%, rgb(239, 239, 239)), linear-gradient(45deg, rgb(239, 239, 239) 25%, transparent 25%, transparent 75%, rgb(239, 239, 239) 75%, rgb(239, 239, 239)); background-position: 0px 0px, 10px 10px; background-size: 21px 21px; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; user-select: none; -webkit-user-drag: none; }

.ndfHFb-c4YZDc-HiaYvf-s2gQvd { inset: 0px; overflow: auto; position: absolute; }

.ndfHFb-c4YZDc-HiaYvf-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { right: initial; }

.ndfHFb-c4YZDc-HiaYvf-haAclf .ndfHFb-c4YZDc-TvD9Pc-qnnXGd, .ndfHFb-c4YZDc-HiaYvf-RJLb9c { height: 100%; position: absolute; width: 100%; }

.ndfHFb-c4YZDc-HiaYvf.ndfHFb-c4YZDc-HiaYvf-gvZm2b-qnnXGd { cursor: crosshair; }

.ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd { box-shadow: rgba(0, 0, 0, 0.5) 0px 2px 4px 0px; border-radius: 3px; position: absolute; z-index: 1; }

.ndfHFb-c4YZDc-HiaYvf-gvZm2b { box-shadow: rgba(0, 0, 0, 0.5) 0px 2px 4px 0px; border-radius: 3px; position: absolute; }

.ndfHFb-c4YZDc-HiaYvf-AHUcCb-oYxtQd.ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd, .ndfHFb-c4YZDc-HiaYvf-gvZm2b { z-index: 2; }

.ndfHFb-c4YZDc-HiaYvf-gvZm2b-SmKAyb, .ndfHFb-c4YZDc-HiaYvf-gvZm2b-n0tgWb { inset: 0px; position: absolute; }

.ndfHFb-c4YZDc-HiaYvf-gvZm2b-SmKAyb { border-radius: 2px; border: 2px solid rgb(255, 255, 255); margin: 1px; z-index: 1; }

.ndfHFb-c4YZDc-HiaYvf-gvZm2b-n0tgWb { border-radius: 3px; border: 2px solid rgba(243, 179, 0, 0.5); z-index: 2; }

.ndfHFb-c4YZDc-HiaYvf-mvZqyf { width: 100%; height: 100%; position: absolute; border: 30000px solid rgb(0, 0, 0); border-radius: 30003px; transform: translate(-30000px, -30000px); opacity: 0; transition: opacity 0.4s ease 0s; pointer-events: none; }

.ndfHFb-c4YZDc-HiaYvf-AHUcCb-oYxtQd .ndfHFb-c4YZDc-HiaYvf-mvZqyf, .ndfHFb-c4YZDc-HiaYvf-gvZm2b .ndfHFb-c4YZDc-HiaYvf-mvZqyf { opacity: 0.5; }

.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd { display: none; }

.ndfHFb-c4YZDc-dkyuHd-ostUZ { position: absolute; min-width: 400px; max-width: 568px; line-height: 20px; top: 8px; background: rgb(26, 115, 232); color: white; overflow: hidden; border-radius: 2px; transform: translate(-50%, -64px); display: flex; align-items: center; box-shadow: rgba(0, 0, 0, 0.5) 0px 2px 4px; transition: transform 0.15s ease 0s; z-index: 4; left: 50%; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ { background: rgb(124, 172, 248); border-radius: 8px; min-width: 364px; box-shadow: none; color: rgb(0, 0, 0); font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); justify-content: space-between; }

.ndfHFb-c4YZDc-dkyuHd-ostUZ.ndfHFb-c4YZDc-dkyuHd-ostUZ-TSZdd { height: auto; transform: translate(-50%, 0px); }

.ndfHFb-c4YZDc-dkyuHd-ostUZ-Ne3sFf { padding: 10px 32px 10px 16px; font-size: 14px; font-weight: 500; float: left; }

.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S, .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:visited { margin-left: auto; margin-top: auto; margin-bottom: auto; text-transform: uppercase; font-size: 14px; cursor: pointer; padding: 10px 16px; text-decoration: none; float: right; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:visited { text-transform: none; width: 24px; height: 24px; }

.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S.ndfHFb-c4YZDc-LgbsSe-XpnDCe, .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:hover { outline: white auto 5px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S .ndfHFb-c4YZDc-Bz112c { background-position: 0px -3570px; width: 24px; height: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S.ndfHFb-c4YZDc-LgbsSe-XpnDCe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:hover { outline: none; }

.ndfHFb-c4YZDc-oKVyEf-haAclf, .ndfHFb-c4YZDc-oKVyEf-haAclf .ndfHFb-c4YZDc-TvD9Pc-qnnXGd { height: 100%; position: absolute; width: 100%; }

.ndfHFb-c4YZDc-oKVyEf-s2gQvd { inset: 0px; overflow: auto; position: absolute; }

.ndfHFb-c4YZDc-oKVyEf-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { right: initial; }

@media print {
  .ndfHFb-c4YZDc-oKVyEf-PEFSMe-OWB6Me { display: none; }
}

.ndfHFb-c4YZDc-SjW3R-ORHb-haAclf { display: none; }

.ndfHFb-c4YZDc-SjW3R-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-SjW3R-ORHb { align-items: center; background: rgb(232, 240, 254); color: rgb(32, 33, 36); display: flex; font-family: "Google Sans", Roboto, arial, sans-serif; height: 48px; width: 100%; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb { background: rgb(124, 172, 248); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-SjW3R-ORHb-haAclf.ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce, .ndfHFb-c4YZDc-SjW3R-ORHb-c6xFrd.ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce, .ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce { display: none; }

.ndfHFb-c4YZDc-SjW3R-ORHb-c6xFrd { align-items: center; display: flex; -webkit-box-flex: 1; flex-grow: 1; float: right; justify-content: flex-end; }

.ndfHFb-c4YZDc-SjW3R-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -2722px; height: 24px; margin: 0px 16px; width: 24px; }

.ndfHFb-c4YZDc-SjW3R-ORHb-Ne3sFf { margin-left: 16px; font-size: 14px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-Bz112c { background-position: 0px -1160px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-Bz112c { background-position: 0px -3570px; }

.ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-sM5MNb { margin: 0px 16px; }

.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover, .ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe { margin: 0px 12px; text-align: center; min-width: 70px; background: rgb(26, 115, 232); border-radius: 5px; font-size: 14px; font-weight: 500; padding: 7px 0px; color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover { background: rgb(43, 125, 233); }

.ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe { margin: 0px 5px; text-align: center; min-width: 70px; color: rgb(26, 115, 232); font-size: 14px; font-weight: 500; padding: 7px 0px; }

.ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover { background: rgb(248, 251, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover { background: transparent; color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-LzGo7c { display: inline-block; font-size: 12px; margin-bottom: 10px; margin-left: 5px; opacity: 0.7; }

.ndfHFb-c4YZDc-LzGo7c-fmcmS { color: rgb(255, 255, 255); display: inline-block; margin-right: 4px; }

.ndfHFb-c4YZDc-LzGo7c .ndfHFb-c4YZDc-LzGo7c-dZ8yzd:link, .ndfHFb-c4YZDc-LzGo7c .ndfHFb-c4YZDc-LzGo7c-dZ8yzd:visited { color: rgb(255, 255, 255); cursor: pointer; display: inline-block; text-decoration: underline; }

.ndfHFb-c4YZDc-hSRGPd-LgbsSe { color: rgb(179, 179, 179); cursor: pointer; text-decoration: underline; }

.ndfHFb-c4YZDc-xl07Ob, .ndfHFb-c4YZDc-mg9Pef { box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; background: rgb(255, 255, 255); color: rgb(51, 51, 51); font-family: arial, sans-serif; font-size: 13px; border: 1px solid rgb(145, 145, 145); line-height: 18px; overflow-y: auto; position: absolute; z-index: 200; outline: transparent solid 1px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob, .ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-mg9Pef { box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 8px; font-family: "Google Sans", Roboto, arial, sans-serif; border: 0px; border-radius: 2px; line-height: 34px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-mg9Pef { background: var(--dt-surface,#fff); border-radius: 4px; }

.ndfHFb-c4YZDc-j7LFlb { cursor: pointer; list-style: none; padding: 6px 6em 6px 37px; position: relative; white-space: nowrap; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb { padding: 1px 60px 1px 52px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb { padding-top: 0px; padding-bottom: 0px; height: 34px; display: flex; align-items: center; }

.ndfHFb-c4YZDc-j7LFlb-Bz112c { background-size: contain; height: 16px; left: 10px; position: absolute; top: 6px; width: 16px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c { left: 16px; height: 20px; width: 20px; }

.ndfHFb-c4YZDc-j7LFlb-sn54Q { background-color: rgb(241, 241, 241); border-color: rgb(241, 241, 241); border-style: dotted; border-width: 1px 0px; padding: 5px 6em 5px 37px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-sn54Q { background-color: rgb(223, 223, 223); border-color: rgb(223, 223, 223); padding: 0px 60px 0px 52px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-sn54Q { background: rgb(55, 55, 55); border: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:hover { background: rgb(47, 47, 47); border: none; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:focus, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:active { background: rgb(55, 55, 55); border: none; }

.ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c { top: 5px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c { top: 6px; }

.ndfHFb-c4YZDc-xl07Ob-tJHJj { color: rgb(89, 89, 89); cursor: default; font-size: 12px; list-style: none; padding: 6px 6em 6px 6px; position: relative; white-space: nowrap; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-tJHJj { padding: 0px 24px 0px 12px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-tJHJj { color: var(--dt-on-surface,#3c4043); }

.ndfHFb-c4YZDc-xl07Ob-hgDUwe { border-bottom: 1px solid rgb(68, 68, 68); }

.ndfHFb-c4YZDc-xl07Ob-WfNeFe-tJHJj { background-color: rgb(239, 239, 239); font-style: italic; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-hgDUwe { border-color: rgb(223, 223, 223); margin: 8px 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-hgDUwe { border-color: var(--dt-outline-variant,#dadce0); margin: 8px 0px; }

.ndfHFb-c4YZDc-mg9Pef .ndfHFb-c4YZDc-j7LFlb { line-height: 36px; padding: 0px 40px 0px 16px; }

.ndfHFb-c4YZDc-mg9Pef .ndfHFb-c4YZDc-j7LFlb-sn54Q { border: none; color: rgba(0, 0, 0, 0.7); }

.ndfHFb-c4YZDc-mg9Pef { padding: 8px 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-bN97Pc { color: var(--dt-on-surface,#3c4043); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-bN97Pc .ndfHFb-c4YZDc-Bz112c { transform: scale(0.83); }

.ndfHFb-c4YZDc-EglORb-haAclf { background-color: rgb(76, 73, 76); border-radius: 12px; color: rgb(255, 255, 255); margin-bottom: 40px; padding: 20px; text-align: center; box-shadow: rgba(0, 0, 0, 0.2) 0px 10px 12px 5px; }

.ndfHFb-c4YZDc-EglORb-haAclf .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c { margin: 0px auto; transform: scale(1.7); }

.ndfHFb-c4YZDc-EglORb-u0pjoe, .ndfHFb-c4YZDc-EglORb-ge6pde, .ndfHFb-c4YZDc-EglORb-Ujd07d { min-width: 300px; position: absolute; text-align: center; }

.ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c { background-repeat: no-repeat; display: inline-block; height: 19px; position: relative; top: 3px; width: 19px; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-spinner_dark.gif") !important; }

.ndfHFb-c4YZDc-e1YmVc.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-spinner_gray.gif") !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { height: 21px; width: 21px; top: 2px; background-image: none !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c .ndfHFb-aZ2wEe { display: block; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c .ndfHFb-vyDMJf-aZ2wEe { height: 32px; width: 32px; margin-left: -16px; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { height: 32px; width: 32px; }

.ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS { font-size: 19px; line-height: 19px; margin-left: 12px; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS { color: rgb(30, 30, 30); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS, .ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS { display: none; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c { background-repeat: no-repeat; background-position: 0px -800px; display: inline-block; height: 37px; margin: 0px auto; padding: 0px; width: 31px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c { background-position: 0px -2424px; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-fmcmS, .ndfHFb-c4YZDc-EglORb-Ujd07d-fmcmS, .ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf { display: inline-block; font-size: 19px; line-height: 27px; user-select: text; }

.ndfHFb-c4YZDc-EglORb-Ujd07d-fmcmS { margin-top: 15px; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf .ndfHFb-c4YZDc-EglORb-u0pjoe-KY1xSc-z5C9Gb-hSRGPd:link, .ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf .ndfHFb-c4YZDc-EglORb-u0pjoe-KY1xSc-z5C9Gb-hSRGPd:visited { padding-left: 5px; color: rgb(255, 255, 255); cursor: pointer; display: inline-block; text-decoration: underline; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb-fmcmS { display: block; font-size: 17px; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb { display: block; font-size: 12px; text-align: left; white-space: pre-wrap; user-select: text; }

.ndfHFb-c4YZDc-EglORb-joDrKf-u0pjoe-fmcmS { font-size: 13px; margin-top: 10px; }

.ndfHFb-c4YZDc-EglORb-u0pjoe-Hr33Cd { font-size: 19px; line-height: 27px; }

.ndfHFb-c4YZDc-EglORb-nupQLb-LgbsSe, .ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe { display: inline-block; }

.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe { margin-left: 20px; margin-top: 20px; border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); font-size: 11px; font-weight: bold; height: 28px; line-height: 28px; min-width: 72px; outline: 0px; padding: 0px 8px; vertical-align: middle; }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.ndfHFb-c4YZDc-LgbsSe-auswjd.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe { background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.ndfHFb-c4YZDc-LgbsSe-XpnDCe.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe { border: 1px solid rgb(77, 144, 254); }

.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-Bz112c { background-size: contain; height: 16px; left: 10px; position: absolute; top: 6px; width: 16px; }

.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-fmcmS { margin-left: 35px; }

.ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf { color: rgb(255, 255, 255); padding-bottom: 20px; text-align: center; }

.ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS { display: inline-block; font-size: 15px; padding-left: 20px; text-align: left; vertical-align: top; }

.XkWAb-LmsqOc, .XkWAb-JaavZc { image-rendering: -webkit-optimize-contrast; }

.XkWAb-LmsqOc { transition: opacity 0.5s linear 0s; }

.XkWAb-xzdHvd { transform: translate(-50%, -50%) rotate(90deg) translate(50%, -50%); }

.XkWAb-hTN0Jd { transform: translate(-50%, -50%) rotate(180deg) translate(-50%, -50%); }

.XkWAb-IZxJAe { transform: translate(-50%, -50%) rotate(270deg) translate(-50%, 50%); }

.XkWAb-cYRDff img.XkWAb-Iak2Lc { transition: none 0s ease 0s; }

.XkWAb-cYRDff img.L6cTce { opacity: 0; }

.XkWAb-CHX6zb { opacity: 0; position: absolute; z-index: 1002; height: 100%; width: 100%; background-color: rgb(0, 128, 0); -webkit-tap-highlight-color: rgba(0, 0, 0, 0); }

.XkWAb-pfZwlb { overflow: hidden; }

.XkWAb-cYRDff { position: absolute; overflow: hidden; background: transparent !important; }

.XkWAb-LmsqOc, .XkWAb-JaavZc { position: absolute; }

.XkWAb-pVNTue { position: absolute; z-index: 1003; width: 1px; height: 1px; user-select: none; }

.XkWAb-RCfa3e { transition: all 0.5s ease 0s; }

.XkWAb-pVNTue.XkWAb-RCfa3e { transition: opacity 0.5s ease 0s; }

.XkWAb-pVNTue .XkWAb-sM5MNb { width: 100%; height: 100%; border: 1px solid rgb(128, 128, 128); background: rgb(0, 0, 0); }

.XkWAb-pVNTue .XkWAb-SMWX4b { direction: ltr; width: 100%; height: 100%; background-repeat: no-repeat; overflow: hidden; position: relative; }

.XkWAb-pVNTue .XkWAb-SMWX4b .XkWAb-pfZwlb .XkWAb-cYRDff { position: absolute; }

.XkWAb-pVNTue .XkWAb-xJ5Hz { border: 1px solid rgb(255, 255, 255); position: absolute; z-index: 1001; background: transparent !important; }

.XkWAb-pVNTue .XkWAb-ZdFRdf { position: absolute; background: rgb(0, 0, 0); opacity: 0.6; z-index: 1001; }

.XkWAb-pVNTue .XkWAb-UH1Jve { width: 100%; height: 30px; background: rgb(0, 0, 0); border-style: solid; border-color: rgb(128, 128, 128); border-width: 0px 1px 1px; position: absolute; transition: height 0.5s ease 0s; }

.XkWAb-eJuzjc, .XkWAb-a4WLyb { color: rgb(255, 255, 255); cursor: pointer; font-size: 13px; height: 30px; position: absolute; top: 0px; text-align: center; transition: height 0.5s ease 0s; vertical-align: middle; width: 22px; }

.XkWAb-BtWyge { display: table-cell; width: 22px; height: 30px; text-align: center; vertical-align: middle; }

.XkWAb-pVNTue .XkWAb-eJuzjc { right: 0px; }

.XkWAb-pVNTue .XkWAb-a4WLyb { left: 0px; }

.XkWAb-pVNTue .XkWAb-IlRY5e { height: 30px; width: 16px; cursor: pointer; transition: height 0.5s ease 0s; background: rgb(255, 255, 255) !important; }

.XkWAb-pVNTue .XkWAb-IE9qgd { left: 22px; position: absolute; right: 22px; top: 0px; transition: height 0.5s ease 0s; }

.XkWAb-AHe6Kc { background-image: url("data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAACAAAAAgAQMAAABJtOi3AAAAAXNSR0IArs4c6QAAAAZQTFRF9/f3////TOsULwAAABRJREFUCNdjYGD4/5+BigR1TWMAAO29P8H0ss2LAAAAAElFTkSuQmCC"); position: absolute; z-index: 1; }

.ndfHFb-c4YZDc-ls4dqb { position: absolute; inset: 0px; z-index: 1; }

.XkWAb-cYRDff, .XkWAb-xJ5Hz { background-color: transparent !important; }

.XkWAb-pVNTue .XkWAb-IlRY5e { background-color: rgb(255, 255, 255) !important; }

.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { opacity: 0.87; background-position: 0px -160px; margin-left: auto; margin-right: auto; margin-top: 3px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-z5C9Gb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-z5C9Gb-LgbsSe-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -400px; margin-top: 2px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-z5C9Gb-LgbsSe-ndfHFb-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1920px; margin-top: 2px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -2746px; margin-top: 0px; height: 24px; width: 24px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1568px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe-ndfHFb-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -328px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-z5C9Gb-xl07Ob { font-size: 13px; min-width: 240px; padding: 8px 0px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-Bz112c { opacity: 0.6; left: 12px; top: 6px; margin-left: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c { top: 5px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c { top: 6px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-z5C9Gb-xl07Ob-xl07Ob-ibnC6b-OWB6Me { opacity: 0.6; }

.ndfHFb-c4YZDc-tJiF1e-LgbsSe, .ndfHFb-c4YZDc-E7ORLb-LgbsSe { position: absolute; top: 80px; bottom: 80px; margin-top: auto; margin-bottom: auto; outline: 0px; width: 40px; height: 90px; z-index: 5; }

.ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1960px; }

.ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -840px; }

.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1640px; }

.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -680px; }

.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c:not([onclick]):not(:link):not(:visited), .ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c:not([onclick]):not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-icons4.png") !important; }

.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: -26px -26px; }

.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -248px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -2096px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -248px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -2096px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe { width: 48px; }

.ndfHFb-c4YZDc-DH6Rkf-Bz112c { height: 24px; position: absolute; width: 24px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-Bz112c { height: 24px; width: 24px; }

.ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { height: 30px; width: 40px; background: rgb(0, 0, 0); border-radius: 3px; opacity: 0.8; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { height: 40px; width: 40px; border-radius: 20px; background: rgba(0, 0, 0, 0.75); transition: background 0.2s ease 0s, opacity 0.34s ease 0s, transform 0.34s cubic-bezier(0.4, 0, 0.2, 1) 0s; opacity: 1; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { background: var(--dt-surface,#fff); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc .ndfHFb-c4YZDc-DH6Rkf-Bz112c { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { background: rgb(66, 133, 244); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { background: rgb(105, 107, 106); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-auswjd .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { background: rgb(109, 111, 111); }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { outline: rgb(77, 144, 254) solid 1px; }

.ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc { display: none; }

.ndfHFb-c4YZDc-zsEIvc-b0t70b { background: white; bottom: 0px; position: absolute; right: 0px; top: 0px; width: 320px; z-index: 4; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-zsEIvc-b0t70b { background: transparent; border-radius: 24px; padding: 0px 16px 16px 0px; box-sizing: border-box; width: 344px; }

.ndfHFb-c4YZDc-zsEIvc-L5Fo6c { border: none; height: 100%; width: 100%; z-index: 4; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-zsEIvc-L5Fo6c { border-radius: 24px; }

@media only screen and (max-width: 500px) {
  .ndfHFb-c4YZDc-zsEIvc-b0t70b { width: 100%; }
}

.ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d { display: inline-block; margin-right: 10px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d { border: 1px solid transparent; border-radius: 2px; background: rgba(0, 0, 0, 0.75); margin: 0px; white-space: nowrap; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d { border-radius: 100px; border-color: var(--dt-outline,#80868b); background-color: var(--dt-surface,#fff); }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe.ndfHFb-c4YZDc-Wrql6b-FNFY6c-BP2Omd-qMHh7d, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c.ndfHFb-c4YZDc-Wrql6b-FNFY6c-BP2Omd-qMHh7d { border-bottom-right-radius: 0px; border-right: 0px; border-top-right-radius: 0px; display: inline-block; margin-right: 0px; min-width: 64px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d { font-size: 13px; font-weight: normal; margin: 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d { min-width: 0px; padding: 0px; color: white; height: 30px; margin-left: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d { color: var(--dt-on-surface-variant,#5f6368); height: 36px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c { padding-right: 4px; min-width: 79px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c { padding-left: 8px; padding-right: 8px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c { padding-left: 16px; padding-right: 16px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d { display: inline-block; min-width: 89px; padding: 10px 0px; }

.ndfHFb-c4YZDc-FNFY6c-V67aGc { display: inline-block; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-V67aGc { line-height: 24px; margin-top: 4px; max-width: 200px; overflow: hidden; text-overflow: ellipsis; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-V67aGc { margin-top: 6px; margin-left: 4px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp { border-bottom-left-radius: 0px; border-left: 0px; border-top-left-radius: 0px; min-width: 15px; }

.ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS { display: inline-block; min-width: 59px; padding-left: 4px; padding-right: 6px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS { line-height: 30px; padding-left: 8px; padding-right: 0px; float: left; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS { line-height: 24px; padding-left: 16px; padding-right: 0px; float: left; margin-top: 4px; }

.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS { display: none; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-PlOyMe, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-FNFY6c, .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-qMHh7d { background-color: rgb(35, 35, 35); background-image: -webkit-linear-gradient(top, rgb(51, 51, 51), rgb(34, 34, 34)); }

.ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb, .ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb { display: inline-block; margin: 0px 4px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb { margin: 0px; overflow: hidden; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb { margin-top: 2px; }

.ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo { opacity: 0.8; display: inline-block; margin-bottom: 1px; vertical-align: middle; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo { opacity: 1; border-bottom-right-radius: 2px; border-right: 2px; border-top-right-radius: 2px; margin-bottom: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo { width: 20px; display: flex; justify-content: center; padding-right: 12px; padding-left: 4px; }

.ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c { background-position: 0px -960px; height: 16px; width: 16px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1936px; height: 24px; width: 24px; margin-top: 4px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c { height: 20px; width: 20px; }

.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo { opacity: 1; }

.ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c { background-size: contain; display: inline-block; height: 16px; margin-right: 6px; width: 16px; vertical-align: text-bottom; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c { float: left; height: 24px; width: 24px; margin-top: 4px; margin-left: -4px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c { height: 14px; width: 14px; margin-top: 11px; margin-bottom: 11px; margin-left: 2px; }

.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe { border-left: 1px solid rgba(255, 255, 255, 0.3); display: inline-block; height: 11px; vertical-align: middle; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe { border-color: rgba(255, 255, 255, 0.35); height: 24px; margin-top: 3px; vertical-align: top; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe { border-color: var(--dt-outline,#80868b); height: 36px; width: 1px; margin-top: 0px; }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE ~ .ndfHFb-c4YZDc-Wrql6b-qMHh7d > .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe, .ndfHFb-c4YZDc-LgbsSe-ZmdkE > .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe { opacity: 0; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE ~ .ndfHFb-c4YZDc-Wrql6b-qMHh7d > .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE > .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe { opacity: 1; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf { transition: opacity 0.218s ease 0s; background-color: rgb(0, 0, 0); border-radius: 3px; bottom: 10px; position: absolute; line-height: 25px; padding: 0px 18px; text-align: center; height: 25px; min-width: 56px; z-index: 3; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-auswjd { opacity: 0.7; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-L6cTce { opacity: 0; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-fmcmS { color: rgb(255, 255, 255); font-size: 11px; font-weight: bold; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb { border-right: 1px solid rgba(255, 255, 255, 0.2); display: inline-block; font-size: 13px; line-height: 44px; height: 44px; vertical-align: middle; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); display: flex; align-items: center; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-tJHJj { display: inline-block; margin-left: 12px; vertical-align: middle; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-DARUcf-NnAfwf-tJHJj { margin-left: 16px; }

.ndfHFb-c4YZDc-DARUcf-NnAfwf-cQYSPc, .ndfHFb-c4YZDc-DARUcf-NnAfwf-j4LONd { display: inline-block; text-align: center; vertical-align: middle; width: 48px; }

.ndfHFb-c4YZDc-cYSp0e, .ndfHFb-c4YZDc-cYSp0e-s2gQvd { inset: 0px; position: absolute; }

.ndfHFb-c4YZDc-cYSp0e-Oz6c3e { position: relative; }

.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e { max-width: 800px; margin: 60px auto; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e { margin-top: 56px; margin-bottom: 56px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e { margin-top: 64px; margin-bottom: 64px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-TJEFFc.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e { margin-top: 12px; margin-bottom: 12px; }

.ndfHFb-c4YZDc-cYSp0e-hpYHOb { bottom: 0px; position: absolute; top: 0px; }

.ndfHFb-c4YZDc-cYSp0e { outline: none; }

.ndfHFb-c4YZDc-cYSp0e-BIzmGd { border: 1px solid rgb(238, 238, 238); box-shadow: rgba(0, 0, 0, 0.05) 0px 3px 3px; background: rgba(255, 255, 255, 0.95); border-radius: 100%; display: block; opacity: 0; position: absolute; width: 40px; height: 40px; left: 100%; margin-left: -22px; cursor: pointer; transition: opacity 0.25s ease-in-out 0s; z-index: 3; }

.ndfHFb-c4YZDc-cYSp0e-BIzmGd.ndfHFb-c4YZDc-LgbsSe { opacity: 1; }

.ndfHFb-c4YZDc-cYSp0e-BIzmGd.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me { opacity: 0; }

.ndfHFb-c4YZDc-BIzmGd-Bz112c { background-position: 0px -2642px; display: inline-block; height: 24px; margin: 10px; opacity: 0.5; pointer-events: none; width: 24px; }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-cYSp0e-BIzmGd .ndfHFb-c4YZDc-BIzmGd-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-cYSp0e-s2gQvd { overflow: auto; }

.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-s2gQvd { margin-left: 12px; margin-right: 12px; overflow: hidden; }

.ndfHFb-c4YZDc-cYSp0e-B7I4Od { left: -5000px; position: absolute; top: -5000px; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf { position: relative; pointer-events: none; background-color: rgba(79, 79, 79, 0.2); }

.ndfHFb-c4YZDc-cYSp0e-DARUcf + .ndfHFb-c4YZDc-cYSp0e-DARUcf { margin-top: 40px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cYSp0e-DARUcf + .ndfHFb-c4YZDc-cYSp0e-DARUcf { margin-top: 16px; }

.ndfHFb-c4YZDc.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-cYSp0e-DARUcf + .ndfHFb-c4YZDc-cYSp0e-DARUcf { margin-top: 12px; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf { font-size: 11px; opacity: 0.01; overflow: hidden; height: 100%; position: absolute; width: 100%; z-index: -1; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj, .ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe { position: absolute; margin: 0px; padding: 0px; border-width: 0px; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-gSKZZ .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf { cursor: text; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-xUXeUb .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf { cursor: crosshair; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c { position: absolute; width: 100%; height: 100%; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-M1R4Ee-UzWXSb { position: absolute; width: 100%; height: 100%; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; background-color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c { box-shadow: none; }

.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf { background-color: transparent; }

.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c { position: relative; height: auto; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf { height: 100%; overflow: hidden; position: absolute; width: 100%; pointer-events: auto; z-index: 2; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-hSRGPd { cursor: pointer; position: absolute; background-image: url("data:image/gif;base64,R0lGODlhAQABAIAAAP///wAAACH5BAEAAAAALAAAAAABAAEAAAICRAEAOw=="); }

.ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q { position: absolute; opacity: 0.35; background-color: rgb(255, 225, 104); z-index: 1; }

.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf, .ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-EglORb-ge6pde { position: relative; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-u0pjoe-DARUcf { position: absolute; height: 100%; width: 100%; pointer-events: auto; z-index: 2; }

.ndfHFb-c4YZDc-cYSp0e-DARUcf-u0pjoe-EglORb { text-align: center; width: 100%; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS { font-size: 15px; line-height: 25px; }

.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c { margin: 5px 0px; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf:not([onclick]):not(:link):not(:visited) { background-color: transparent !important; }

.ndfHFb-c4YZDc-UmsTj-Sx9Kwc { position: absolute; min-width: 400px; height: 105px; background: rgb(35, 35, 35); border: 1px solid rgb(0, 0, 0); border-radius: 3px; color: white; cursor: default; font-size: 15px; font-weight: bold; font-family: arial, sans-serif; user-select: text; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc { background: var(--dt-surface,#fff); padding: 24px; border-radius: 8px; display: flex; align-items: center; flex-direction: column; justify-content: space-between; height: auto; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc-ma6Yeb { display: flex; flex-direction: row; margin: 0px 0px 24px; }

.ndfHFb-c4YZDc-UmsTj-Ne3sFf { position: relative; top: 11px; margin-left: 40px; margin-right: 10px; white-space: nowrap; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Ne3sFf { position: static; font: var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-large-spacing,0); margin: 0px 16px; }

.ndfHFb-c4YZDc-UmsTj-Bz112c { position: absolute; top: 4px; left: 7px; width: 28px; height: 28px; background-position: 0px -920px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UmsTj-Bz112c { background-position: 0px -1328px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UmsTj-Bz112c { background-position: 0px -472px; position: static; }

.ndfHFb-c4YZDc-UmsTj-YPqjbf-sM5MNb { position: absolute; left: 10px; right: 10px; top: 40px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-YPqjbf-sM5MNb { position: static; width: 100%; }

.ndfHFb-c4YZDc-UmsTj-YPqjbf { position: absolute; top: 0px; height: 19px; width: 100%; margin: 0px; background-color: rgb(92, 92, 92); border: 1px solid rgb(0, 0, 0); color: white; font: 16px arial, sans-serif; box-sizing: content-box; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-YPqjbf { position: static; height: 26px; box-sizing: border-box; }

.ndfHFb-c4YZDc-UmsTj-Sx9Kwc-cGMI2b { position: relative; top: 53px; width: 100%; white-space: nowrap; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc-cGMI2b { position: static; display: flex; flex-direction: row; justify-content: space-between; margin: 24px 0px 0px; }

.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf { top: 0px; right: 9px; background-color: rgb(77, 144, 254); color: rgba(255, 255, 255, 0.87); margin: 0px; padding: 0px 8px; font-size: 13px; height: 25px; line-height: 25px; min-width: 50px; text-align: center; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf { border-radius: 100px; background: var(--dt-surface,#fff); color: var(--dt-primary,#1a73e8); font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; font-size: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); border: none; margin: 0px; padding: 0px; position: static; height: 30px; min-width: 72px; line-height: 30px; }

.ndfHFb-c4YZDc-UmsTj-u0pjoe { top: 2px; min-width: 295px; white-space: nowrap; display: inline-block; position: static; margin: 0px; }

.ndfHFb-c4YZDc-UmsTj-u0pjoe-fmcmS { color: rgb(255, 0, 0); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-u0pjoe-fmcmS { color: var(--dt-error,#d93025); font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; font-size: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-large-spacing,0.00625em); height: 30px; line-height: 30px; }

.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-UmsTj-sFeBqf { background-color: rgb(128, 128, 128); color: rgb(194, 194, 194); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-UmsTj-sFeBqf { background: var(--dt-surface,#fff); color: var(--dt-on-surface,#3c4043); opacity: 0.38; }

.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-UmsTj-sFeBqf { background-color: rgb(77, 144, 254); background-image: -webkit-linear-gradient(top, rgb(77, 144, 254), rgb(53, 122, 232)); color: rgb(255, 255, 255); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-UmsTj-sFeBqf { background: rgba(168, 199, 250, 0.08); color: var(--dt-primary,#1a73e8); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf:active { background: rgba(168, 199, 250, 0.12); color: var(--dt-primary,#1a73e8); border: none; outline: none; box-shadow: none; }

.ndfHFb-c4YZDc-ujibv-nUpftc { display: block; margin-left: 12px; margin-right: 12px; margin-top: 56px; z-index: 1; }

.ndfHFb-c4YZDc-ujibv-nUpftc .ndfHFb-c4YZDc-ujibv-JUCs7e { left: 50%; max-width: max-content; position: relative; transform: translateX(-50%); width: 100%; }

.ndfHFb-c4YZDc-n1UuX-Bz112c, .ndfHFb-c4YZDc-mKZypf-bEDTcc, .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-yHKmmc, .ndfHFb-c4YZDc-no16zc-UcSZ6e { display: inline-block; padding: 9px 0px; }

.ndfHFb-c4YZDc-Woal0c-jcJzye-ZMv3u { vertical-align: middle; }

.ndfHFb-c4YZDc-n1UuX-RJLb9c { background-color: rgb(70, 68, 69); border-radius: 50%; height: 29px; width: 29px; margin-left: 13px; vertical-align: middle; }

.ndfHFb-c4YZDc-no16zc-UcSZ6e { vertical-align: middle; }

.ndfHFb-c4YZDc-no16zc-UcSZ6e-LgbsSe { margin-left: 13px; margin-right: 0px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.ndfHFb-c4YZDc-mKZypf-bEDTcc-LgbsSe { margin-left: 13px; margin-right: 0px; }

.ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe, .ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe { display: inline-block; margin-left: 13px; margin-right: 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-n1UuX-Bz112c { padding: 5.5px 8px; margin-left: 3px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-mKZypf-bEDTcc, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-yHKmmc, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-no16zc-UcSZ6e { padding: 5.5px 8px; margin-left: 8px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-n1UuX-RJLb9c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-mKZypf-bEDTcc-LgbsSe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-no16zc-UcSZ6e-LgbsSe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe { margin-left: 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe + .ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe { margin-left: 13px; }

.ndfHFb-c4YZDc-kODWGd-umzg3c { height: 100%; position: absolute; left: 46px; right: auto; }

.ndfHFb-c4YZDc-kODWGd-umzg3c-SxecR { width: 130px; }

.ndfHFb-c4YZDc-kODWGd-umzg3c-SxecR-PFprWc { height: 12px; width: 20px; }

.ndfHFb-c4YZDc-kODWGd-umzg3c-ihIZgd { font-family: "Open Sans", arial, sans-serif; font-size: 13px; font-weight: bold; min-width: 30px; top: 8px; left: 144px; right: auto; position: absolute; }

.ndfHFb-c4YZDc-sbW6Cb { box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; background-color: rgb(248, 248, 248); color: rgb(42, 42, 42); display: block; font: 13px / 19px "Google Sans", arial, sans-serif; margin-left: 20px; opacity: 1; position: absolute; visibility: visible; z-index: 201; }

.ndfHFb-c4YZDc-sbW6Cb-bN97Pc { padding: 10px; }

.ndfHFb-c4YZDc-sbW6Cb-bN97Pc-hSRGPd { color: rgb(42, 42, 42); text-decoration: underline; }

.ndfHFb-c4YZDc-sbW6Cb-hFsbo { position: absolute; }

.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe, .ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { content: ""; display: block; height: 0px; position: absolute; width: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe { border: 16px solid; }

.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border: 14px solid; }

.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb { bottom: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-d6mlqf { top: -14px; }

.ndfHFb-c4YZDc-sbW6Cb-y6n2Me { left: -14px; }

.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc { right: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe, .ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe { border-color: rgb(248, 248, 248) transparent; left: -16px; }

.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc, .ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-color: rgb(248, 248, 248) transparent; left: -14px; }

.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe, .ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-bottom-width: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe { border-top-width: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-top-width: 0px; top: 2px; }

.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe, .ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe { border-color: transparent rgb(248, 248, 248); top: -16px; }

.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc, .ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-color: transparent rgb(248, 248, 248); top: -14px; }

.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe { border-left-width: 0px; }

.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-left-width: 0px; left: 2px; }

.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe, .ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc { border-right-width: 0px; }

.ndfHFb-c4YZDc-Lo93Wb-fmcmS { display: inline-block; vertical-align: middle; max-width: 150px; margin-right: 5px; }

.ndfHFb-c4YZDc-Lo93Wb-Bz112c { display: inline-block; vertical-align: middle; background-repeat: no-repeat; opacity: 0.87; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc { color: rgb(0, 0, 0); font: 13px arial, sans-serif; width: 340px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc { color: var(--dt-on-surface,#3c4043); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-r4nke { font-weight: normal; margin: 0px 0px 16px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-r4nke { margin: 0px 0px 24px; }

.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc { border-radius: 1px; border-width: 1px; border-style: solid; border-color: rgb(192, 192, 192) rgb(217, 217, 217) rgb(217, 217, 217); border-image: initial; font-size: 13px; height: 25px; padding: 1px 8px; width: 300px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc { border: 2px solid var(--dt-primary,#1a73e8); font: var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-large-spacing,0.00625em); padding: 8px 16px; border-radius: 4px; background: var(--dt-surface,#fff); color: var(--dt-on-surface,#3c4043); }

.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc:focus { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; border: 1px solid rgb(77, 144, 254); outline: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc:focus { border: 2px solid var(--dt-primary,#1a73e8); }

.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd { margin-top: 16px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd { margin-top: 24px; display: flex; justify-content: flex-end; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd button { cursor: pointer; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Iqlsrf-Bz112c { background-position: 0px -976px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Iqlsrf-Bz112c { background-position: 0px -856px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-bN97Pc br { display: none; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe { position: absolute; left: -300px; top: -42px; z-index: 4; height: 40px; width: 295px; background-color: rgb(45, 45, 45); border: 1px solid rgb(0, 0, 0); border-radius: 3px; transition: top 0.218s ease-out 0s; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe { left: -600px; background: var(--dt-surface3,#fff); box-shadow: rgba(0, 0, 0, 0.15) 0px 4px 8px 3px, rgba(0, 0, 0, 0.3) 0px 1px 3px; border-radius: 8px; padding: 12px 16px; border: none; height: 36px; display: flex; align-items: center; width: 336px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-ti6hGc, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-ti6hGc { left: unset; right: 56px; top: 50px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf { position: relative; margin: 0px 0px 0px 4px; vertical-align: middle; height: 25px; padding: 0px 9px; width: 198px; background-color: rgb(10, 10, 10); border-style: solid; border-color: rgb(68, 68, 68); border-image: initial; border-width: 0px 0px 1px 1px; display: inline-block; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf { display: flex; align-items: center; width: 200px; height: auto; margin: 0px; padding: 4px 8px; background: var(--dt-surface3,#fff); border: 1px solid var(--dt-outline,#80868b); border-radius: 4px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf:hover { border: 1px solid var(--dt-on-surface,#3c4043); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf-XpnDCe { border: 2px solid var(--dt-primary,#1a73e8); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-x5ghY { border: 2px solid var(--dt-error,#d93025); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf-haAclf { display: table-cell; width: 100%; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf, .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf { color: rgb(255, 255, 255); font-size: 13px; font-weight: normal; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf { width: 100%; background-color: rgb(10, 10, 10); border: 0px; height: 25px; padding: 0px; outline: none !important; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf { height: 24px; font: var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-large-spacing,0.00625em); background: var(--dt-surface3,#fff); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf::-webkit-input-placeholder { color: rgb(255, 255, 255); opacity: 0.75; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-haAclf { display: table-cell; max-width: 100px; opacity: 0.5; padding-left: 7px; white-space: nowrap; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf { padding: 0px 2px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-x5ghY { background-color: rgb(255, 69, 0); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-y7UsZc { display: inline-block; height: 100%; position: absolute; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne { position: relative; top: 8px; height: 21px; width: 21px; opacity: 0.7; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne { position: static; top: 0px; opacity: 1; border-radius: 100px; margin-left: 8px; padding: 8px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne { opacity: 0.9; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne { opacity: 1; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgba(196, 199, 197, 0.08); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-XpnDCe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-auswjd { background-color: rgba(196, 199, 197, 0.12); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc { background-position: 0px 0px; margin-left: -2px; top: 5px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc { top: 0px; margin-left: 8px; height: 21px; width: 21px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc .ndfHFb-c4YZDc-Bz112c { transform: scale(0.86); position: relative; top: -1px; right: 1px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc.ndfHFb-c4YZDc-w5vlXd { top: 8px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc.ndfHFb-c4YZDc-w5vlXd { top: -1px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e, .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb { border: 1px solid rgb(68, 68, 68); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb { border: none; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e { background-position: 0px -80px; left: -1px; border-top-right-radius: 3px; border-bottom-right-radius: 3px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e .ndfHFb-c4YZDc-Bz112c { position: relative; top: 1px; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb { background-position: 0px -1240px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc { background-position: 0px -3178px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e { background-position: 0px -1752px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb { background-position: 0px -3754px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne .ndfHFb-c4YZDc-Bz112c { height: 21px; width: 21px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc .ndfHFb-c4YZDc-Bz112c { background-position: 0px -3178px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1752px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb .ndfHFb-c4YZDc-Bz112c { background-position: 0px -3754px; }

.ndfHFb-c4YZDc-O1htCb-LgbsSe, .ndfHFb-c4YZDc-O1htCb-K2kob { background-color: rgba(90, 90, 90, 0.7); border: 2px solid rgb(215, 215, 215); height: 32px; left: 70px; position: absolute; top: 80px; width: 32px; z-index: 5; border-radius: 50%; }

@media screen and (max-width: 800px) {
  .ndfHFb-c4YZDc-O1htCb-LgbsSe { left: 5%; }
}

.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE, .VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-O1htCb-K2kob { background-color: rgba(138, 138, 138, 0.7); border: 2px solid rgb(255, 255, 255); box-shadow: rgba(83, 83, 83, 0.7) 0px 2px 5px; }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe, .VIpgJd-wQNmvb-gk6SMd .ndfHFb-c4YZDc-O1htCb-K2kob { background-color: rgb(77, 144, 254); border: 2px solid rgb(255, 255, 255); box-shadow: rgba(83, 83, 83, 0.7) 0px 2px 5px; }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE, .VIpgJd-wQNmvb-gk6SMd.VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-O1htCb-K2kob { background-color: rgb(94, 155, 254); }

.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-O1htCb-LgbsSe-gk6SMd-YLEHIf, .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b-YLEHIf .ndfHFb-c4YZDc-O1htCb-K2kob { animation: 0.3s linear 0s 1 normal none running driveViewerSelectButtonSelectedAnimation; }

.ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c, .ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg"); background-position: 0px -1320px; width: 30px; height: 30px; margin-top: -4px; opacity: 0.7; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c, .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -2682px; }

.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c { opacity: 0.9; }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c { opacity: 1; }

@-webkit-keyframes driveViewerSelectButtonSelectedAnimation { 
  0% { opacity: 0.3; transform: scale(0.7); }
  50% { opacity: 1; transform: scale(1.1); }
  70% { transform: scale(0.9); }
  100% { transform: scale(1); }
}

@keyframes driveViewerSelectButtonSelectedAnimation { 
  0% { opacity: 0.3; transform: scale(0.7); }
  50% { opacity: 1; transform: scale(1.1); }
  70% { transform: scale(0.9); }
  100% { transform: scale(1); }
}

.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob { background: rgb(237, 237, 237); border-radius: 3px; border: none; box-shadow: rgba(0, 0, 0, 0.4) 0px 1px 2px 1px; margin-top: 4px; margin-left: -35px; max-height: 70%; max-width: 645px; }

.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-j7LFlb { display: inline-block; padding: 0px; }

.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q { padding: 0px; border: none; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-JUCs7e { border: none; border-radius: 0px; display: block; height: auto; margin: 0px; width: auto; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b { display: inline-block; height: 110px; margin: 3px 8px; overflow: hidden; position: relative; width: 110px; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-JUCs7e-SmKAyb { display: table-cell; height: 90px; text-align: center; vertical-align: middle; width: 110px; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-JUCs7e-SmKAyb img { box-shadow: rgba(0, 0, 0, 0.7) 0px 1px 2px 0px; max-width: 100%; max-height: 90%; display: inline-block; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b img.ndfHFb-c4YZDc-JUCs7e-Bz112c { background-color: rgb(245, 245, 245); height: 60px; width: 60px; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b-r4nke { font-size: 15px; margin-top: 3px; overflow: hidden; text-overflow: ellipsis; text-align: center; white-space: nowrap; }

@media screen and (max-width: 1350px) {
  .ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob { max-width: 520px; }
}

@media screen and (max-width: 1000px) {
  .ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob { max-width: 390px; }
}

@media screen and (max-width: 700px) {
  .ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob { max-width: 273px; }
}

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob { position: absolute; right: 0px; top: 55px; }

.VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob, .VIpgJd-wQNmvb-gk6SMd .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob { box-shadow: none; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-wQNmvb-gk6SMd { background-image: none; }

.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-j7LFlb-sn54Q, .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-j7LFlb-ZmdkE { background-color: transparent; border: none; padding: 0px; }

.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf { padding: 0px; }

.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd { padding: 14px 24px 4px; display: flex; border: none; background: rgb(31, 31, 31); color: rgb(227, 227, 227); height: 30px; }

.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf .euCgFf-PLEiK-hSRGPd { text-transform: none; border-radius: 100px; height: 30px; margin: 0px 0px 0px 16px; padding: 0px 16px; color: rgb(168, 199, 250); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf .euCgFf-PLEiK-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf .euCgFf-PLEiK-Bz112c { margin-right: 8px; }

.ndfHFb-c4YZDc-ZCZpd-h9d3hd { box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; outline: none; z-index: 200 !important; }

.ndfHFb-c4YZDc-qbOKL-OEVmcd .IyROMc-w3KqTd-ztA2jd-SUR3Rd { z-index: 201 !important; }

.ndfHFb-c4YZDc-SxecR { height: 12px; margin-top: 12px; padding-left: 0px; padding-right: 2px; }

.ndfHFb-c4YZDc-SxecR-PFprWc { background-image: -webkit-linear-gradient(top, rgb(255, 255, 255), rgb(192, 192, 192)); box-shadow: rgb(0, 0, 0) 0px 0px 5px 0px; border-radius: 6px; position: absolute; top: 10px; background-color: rgb(229, 229, 229) !important; }

.ndfHFb-c4YZDc-SxecR-skjTt { border-radius: 8px; height: 6px; position: absolute; }

.ndfHFb-c4YZDc-SxecR-cQwEuf { background-color: rgb(77, 77, 77); margin-top: 1px; width: 0px; }

.ndfHFb-c4YZDc-SxecR-skjTt-j4LONd { background-color: transparent; width: inherit; border: 1px solid rgb(128, 128, 128) !important; }

.ndfHFb-c4YZDc-SxecR-skjTt-MFS4be { background-image: -webkit-linear-gradient(top, rgb(195, 195, 195), rgb(217, 217, 217)); border-bottom-right-radius: 0px; border-top-right-radius: 0px; margin-top: 1px; width: 0px; background-color: rgb(217, 217, 217) !important; }

.ndfHFb-c4YZDc-Ng57nc.ndfHFb-c4YZDc-b3rLgd-haAclf { bottom: 24px; left: 24px; position: absolute; text-align: left; z-index: 4; }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc.ndfHFb-c4YZDc-b3rLgd-haAclf { bottom: 0px; left: 0px; text-align: center; width: 100%; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd { border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; align-items: center; display: flex; transform: translate3d(0px, 72px, 0px); transition: transform 0.15s cubic-bezier(0.4, 0, 1, 1) 0s, opacity 0.15s cubic-bezier(0.4, 0, 1, 1) 0s, visibility 0ms linear 0.15s; background-color: rgb(238, 238, 238); border: none; color: black; font-size: 14px; margin: 0px; max-width: 568px; min-height: 20px; min-width: 288px; opacity: 0; padding: 14px 0px 14px 24px; text-align: left; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd { background: var(--dt-surface,#fff); color: var(--dt-on-surface,#3c4043); padding: 14px 8px 14px 24px; }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd { background-color: rgb(50, 50, 50); color: white; max-width: none; width: 100%; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-TSZdd { transition-delay: 0s; transform: translate3d(0px, 0px, 0px); bottom: 24px; opacity: 1; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-Ne3sFf { align-items: center; display: flex; flex: 1 1 0px; line-height: 19px; overflow: hidden; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd { flex: 0 0 auto; padding-left: 24px; padding-right: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd { text-transform: none; border-radius: 100px; height: 30px; line-height: 30px; margin: 0px 8px 0px 16px; padding: 0px 16px; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited { background: none; border: none; color: rgb(25, 103, 210); cursor: pointer; font-family: inherit; font-size: inherit; font-weight: bold; margin: 0px; outline: none; text-decoration: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited { color: var(--dt-primary,#1a73e8); }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited { text-transform: uppercase; float: right; }

.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover, .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:focus { text-decoration: underline; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:focus { text-decoration: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover { background: rgba(168, 199, 250, 0.08); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:active { background: rgba(168, 199, 250, 0.12); }

.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd { color: rgb(161, 194, 250); padding-right: 48px; }

.ndfHFb-c4YZDc-L7w45e-ORHb { display: none; align-items: center; background-color: rgb(249, 171, 0); border-radius: 0px; color: rgb(32, 33, 36); height: 3rem; position: relative; top: 0px; width: 100%; z-index: 3; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb { background: rgb(255, 223, 153); }

.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb { display: none; align-items: center; background-color: var(--dt-error,#d93025); border-radius: 0px; color: rgb(255, 255, 255); height: 3rem; position: relative; top: 0px; width: 100%; z-index: 3; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb { background: rgb(236, 146, 142); color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-L7w45e-ORHb.ndfHFb-c4YZDc-ORHb-ZiwkRe, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb.ndfHFb-c4YZDc-ORHb-ZiwkRe { display: flex; }

.ndfHFb-c4YZDc-L7w45e-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3098px; height: 24px; margin: 0px 25px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Bz112c { margin: 0px 16px; }

.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3714px; height: 24px; margin: 0px 25px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Bz112c { background-position: 0px -3098px; margin: 0px 16px; }

.ndfHFb-c4YZDc-L7w45e-ORHb-bN97Pc, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-bN97Pc { align-items: center; display: flex; justify-content: space-between; width: 100%; }

.ndfHFb-c4YZDc-L7w45e-ORHb-Ne3sFf, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Ne3sFf { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Ne3sFf, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Ne3sFf { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,0.0142857143em); }

.ndfHFb-c4YZDc-L7w45e-ORHb-LQLjdd, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-LQLjdd { display: flex; align-items: center; margin: 8px 0px; order: 0; }

.ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3570px; }

.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c { background-image: url("//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg"); background-position: 0px -3178px; }

.ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-Bz112c, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c { margin: 0px 16px; height: 20px; width: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c { background-position: 0px -3570px; }

.ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe { align-self: center; color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; padding: 4px 18px; text-align: center; text-decoration: none; border-radius: 20px; border: 1px solid black; }

.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe { align-self: center; color: rgb(255, 255, 255); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; padding: 4px 18px; text-align: center; text-decoration: none; border-radius: 20px; border: 1px solid white; }

.ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe { align-self: center; color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; padding: 0px 16px; text-align: center; text-decoration: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe { border: none; color: rgb(32, 33, 36); font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); padding: 0px 12px; min-width: 70px; }

.ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe:hover, .ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe:hover, .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe:hover { cursor: pointer; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc { align-items: flex-start; display: flex; flex-direction: column; padding: 0px; outline: none; position: absolute; width: 468px; background: rgb(255, 255, 255); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; border-radius: 8px; z-index: 101; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc { background: var(--dt-surface,#fff); padding: 24px; border-radius: 8px; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); height: 100%; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 101; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-bN97Pc { color: rgb(241, 243, 244); display: flex; flex-direction: column; justify-content: space-between; margin: 0px 12px 12px; text-align: left; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-bN97Pc { background-color: var(--dt-surface,#fff); margin: 0px; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke { margin: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke { margin: 0px; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1.375rem; font-weight: 400; letter-spacing: 0px; line-height: 1.75rem; color: rgb(32, 33, 36); }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke-fmcmS { background-color: var(--dt-surface,#fff); color: var(--dt-on-surface,#3c4043); font: var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-headline-small-spacing,0); }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-g7W7Ed { color: rgb(32, 33, 36); font-family: Roboto; font-style: normal; font-weight: 400; font-size: 14px; line-height: 20px; letter-spacing: 0.2px; margin-bottom: 22.6px; width: 428px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-g7W7Ed { font: var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-large-spacing,0.00625em); margin: 24px 0px; color: var(--dt-on-surface,#3c4043); }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-c6xFrd { margin-right: 22px; margin-left: auto; margin-bottom: 18px; display: flex; flex-direction: row; padding: 0px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-c6xFrd { margin: 0px; display: flex; flex-direction: row; width: 100%; justify-content: flex-end; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 20px; border: none; background: rgb(26, 115, 232); box-sizing: border-box; border-radius: 4px; color: rgb(255, 255, 255); margin: 0px 12px; min-width: 70px; outline: none; padding: 8px 24px; text-align: center; cursor: pointer; }

.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 14px; line-height: 20px; background: rgb(255, 255, 255); border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(26, 115, 232); margin: 0px 12px; min-width: 70px; outline: none; padding: 8px 24px; text-align: center; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe { margin: 0px 0px 0px 24px; border-radius: 100px; background: var(--dt-surface,#fff); color: var(--dt-primary,#1a73e8); font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,0.0178571429em); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:hover, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:hover { background: rgba(168, 199, 250, 0.08); color: var(--dt-primary,#1a73e8); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:active, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:active { background: rgba(168, 199, 250, 0.12); color: var(--dt-primary,#1a73e8); border: none; outline: none; box-shadow: none; }

.ndfHFb-c4YZDc-Wrql6b { background-color: rgba(0, 0, 0, 0.6); height: 27px; padding: 10px 0px; position: absolute; top: 0px; width: 100%; z-index: 3; }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b { background-color: rgb(77, 144, 254); }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b { background-color: rgba(147, 147, 147, 0.7); padding: 10px 0px; }

.ndfHFb-c4YZDc-Wrql6b-hOcTPc { left: 20px; position: absolute; white-space: nowrap; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Wrql6b-hOcTPc { display: flex; align-items: center; position: static; }

.ndfHFb-c4YZDc-Wrql6b-hOcTPc .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c { float: right; }

.ndfHFb-c4YZDc-Wrql6b-LQLjdd { position: absolute; top: 0px; white-space: nowrap; height: 47px; }

.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd { background-color: rgb(77, 144, 254); border-left: 1px solid rgb(106, 163, 255); border-right: 1px solid rgb(106, 163, 255); }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b-LQLjdd { border-color: transparent; }

.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b { display: inline-block; }

.ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b { position: absolute; right: 16px; top: 0px; white-space: nowrap; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b { right: 0px; }

.ndfHFb-c4YZDc-Wrql6b-N7Eqid { background-color: rgba(0, 0, 0, 0.6); display: inline-block; font-size: 11px; line-height: 28px; margin-right: 10px; vertical-align: top; }

.ndfHFb-c4YZDc-Wrql6b-Bz112c { background-size: contain; display: inline-block; float: left; height: 16px; margin-right: 12px; position: relative; top: 8px; width: 16px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Wrql6b-Bz112c { top: 0px; }

.ndfHFb-c4YZDc-Wrql6b-jfdpUb { color: rgb(179, 179, 179); display: inline-block; }

.ndfHFb-c4YZDc-Wrql6b-V1ur5d { color: rgb(255, 255, 255); font-size: 13px; font-weight: normal; line-height: 27px; }

.ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-qnnXGd { line-height: 20px; }

.ndfHFb-c4YZDc-Wrql6b-V1ur5d-hpYHOb, .ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-hpYHOb { visibility: hidden; position: absolute; height: auto; width: auto; }

.ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Iqlsrf-qnnXGd { cursor: pointer; }

.ndfHFb-c4YZDc-Wrql6b-V1ur5d-hSRGPd:hover { cursor: pointer; text-decoration: underline; }

.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d { font-size: 11px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b { pointer-events: none; background: linear-gradient(rgba(0, 0, 0, 0.65) 0%, transparent 100%); height: 56px; padding: 0px 0px 16px; left: 0px; right: 0px; width: auto; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b { height: 64px; padding: 0px; background: transparent; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b.ndfHFb-c4YZDc-Wrql6b-Hyc8Sd { height: 64px; padding: 0px; background: rgba(31, 31, 31, 0.85); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-SmKAyb { position: absolute; pointer-events: auto; height: 48px; left: 0px; right: 0px; padding-top: 8px; width: auto; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-SmKAyb { display: flex; justify-content: space-between; align-items: center; padding-top: 0px; height: 64px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b.ndfHFb-c4YZDc-Wrql6b-qbOKL { box-shadow: rgba(0, 0, 0, 0.6) 0px 2px 2px; background: rgb(50, 50, 50); padding: 0px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b { background: rgba(0, 0, 0, 0.75); height: 40px; top: 12px; left: auto; padding: 0px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-SmKAyb { height: 40px; padding: 0px; margin: 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { margin-left: 8px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-DdWCyb-b0t70b { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b { top: auto; right: 0px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b { display: flex; position: static; align-items: center; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b.ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b-SfQLQb-Woal0c-jcJzye-n1UuX { top: 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-Bz112c { border-radius: 2px; margin: 3px 11px; width: 18px; height: 18px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-jfdpUb { letter-spacing: 0px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d { font-size: 14px; line-height: 40px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,0.00625em); }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-qnnXGd { line-height: 30px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-LQLjdd { display: inline-block; position: relative; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-LQLjdd { display: flex; align-items: center; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { float: left; margin-left: 0px; }

.ndfHFb-c4YZDc-hDEnYe { width: 100%; height: 100%; padding-top: 47px; box-sizing: border-box; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-hDEnYe { padding-top: 0px; }

.ndfHFb-c4YZDc-i5oIFb:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-hDEnYe { padding-top: 56px; }

.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-hDEnYe { padding-top: 64px; }

.ndfHFb-c4YZDc-hDEnYe-SmKAyb { width: 100%; height: 100%; box-sizing: border-box; padding-bottom: 39px; }

.ndfHFb-c4YZDc-hDEnYe-SmKAyb .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { position: relative; right: initial; top: initial; }

.ndfHFb-c4YZDc-hDEnYe-AznF2e { width: 100%; height: 100%; font-size: 0px; box-sizing: border-box; position: relative; }

.ndfHFb-c4YZDc-hDEnYe-AznF2e > .ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-hDEnYe-XuHpsb-haAclf { background-color: transparent; z-index: 1; overflow: auto; position: absolute; inset: 0px; }

.ndfHFb-c4YZDc-hDEnYe-RwANvf-BvBYQ-haAclf { position: absolute; left: 0px; bottom: 0px; overflow-y: hidden; }

.ndfHFb-c4YZDc-hDEnYe-RwANvf-DKlKme-haAclf { position: absolute; top: 0px; overflow-x: hidden; }

.ndfHFb-c4YZDc-hDEnYe-RwANvf-qbOKL-PLDbbf { position: absolute; overflow: hidden; }

.ndfHFb-c4YZDc-hDEnYe-XuHpsb-qJTHM { position: relative; }

.ndfHFb-c4YZDc-hDEnYe-Df1ZY-bN97Pc { font-size: 11px; opacity: 0.01; overflow: hidden; position: absolute; width: 100%; height: 100%; left: 0px; top: 0px; z-index: -1; display: block; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc { width: 100%; z-index: 3; background-color: rgb(0, 0, 0); position: absolute; bottom: 0px; padding-left: 46px; box-sizing: border-box; white-space: nowrap; padding-bottom: 6px; padding-top: 1px; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { font-size: 12px; font-weight: normal; padding: 0px 8px; max-width: 200px; overflow: hidden; background-color: rgb(33, 33, 33); background-image: none; color: rgb(152, 152, 152); line-height: 32px; margin-right: 4px; border: none; border-radius: 0px 0px 3px 3px; height: inherit; box-shadow: none; text-overflow: ellipsis; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { padding: 5px 0px 1px; }

.ndfHFb-c4YZDc-hDEnYe-z5C9Gb-Bz112c { background-position: 0px -200px; width: 24px; height: 24px; margin-left: auto; margin-right: auto; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hDEnYe-z5C9Gb-Bz112c { background-position: 0px -2056px; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe { background-color: rgb(74, 74, 74); color: white; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { color: white; cursor: pointer; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob { background-color: rgb(33, 33, 33); border: none; max-height: 200px; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob > .ndfHFb-c4YZDc-j7LFlb { margin: 0px 20px; padding: 0px; font-size: 12px; color: rgb(152, 152, 152); height: 32px; border: none; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob > .ndfHFb-c4YZDc-j7LFlb > .ndfHFb-c4YZDc-j7LFlb-bN97Pc { max-width: 250px; min-width: 30px; white-space: nowrap; text-overflow: ellipsis; overflow-x: hidden; line-height: 32px; display: inline-block; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob > .ndfHFb-c4YZDc-j7LFlb-sn54Q { color: white; cursor: pointer; background-color: inherit; }

.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob > .ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-j7LFlb { background-color: rgb(74, 74, 74); color: white; }

.ndfHFb-c4YZDc-hDEnYe-eFD6re { left: -5000px; position: absolute; top: -5000px; }

.ndfHFb-c4YZDc-hDEnYe-wvGCSb-gkA7Yd-haAclf .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { left: 30px; position: absolute; right: 30px; top: 0px; }

.ndfHFb-c4YZDc-hDEnYe-wvGCSb-gkA7Yd-haAclf { inset: 56px 0px 39px auto; overflow: auto; padding-top: 8px; position: absolute; width: 362px; }

.ndfHFb-c4YZDc-hDEnYe-wvGCSb-bF1uUb { inset: 56px 0px 39px; overflow: hidden; position: absolute; }

.ndfHFb-c4YZDc-hDEnYe-jNm5if-Bz112c-awotqb { display: inline-block; margin: 0px 4px; vertical-align: middle; }

.ndfHFb-c4YZDc-hDEnYe-jNm5if-NnAfwf-VCkuzd { background: white; border-radius: 2px 2px 0px; color: black; height: 16px; min-width: 12px; padding: 0px 4px; position: relative; text-align: center; top: -1px; }

.ndfHFb-c4YZDc-hDEnYe-jNm5if-NnAfwf { font-family: "Google Sans", Roboto, arial, sans-serif; font-size: 10px; position: relative; top: -9px; }

.ndfHFb-c4YZDc-hDEnYe-jNm5if-Zj4Smb { border-left: 4px solid transparent; border-top: 4px solid white; height: 0px; position: absolute; right: 0px; top: 16px; width: 0px; }

.ndfHFb-c4YZDc-hDEnYe-wvGCSb-ge6pde-uDEFge { background: rgb(66, 133, 244); left: 50%; padding: 10px 16px; position: absolute; top: 68px; transform: translateX(-50%); }

.ndfHFb-c4YZDc-hDEnYe-XuHpsb-hSRGPd-haAclf { user-select: none; }

.ndfHFb-c4YZDc-hDEnYe-bN97Pc { position: absolute; }

.ndfHFb-c4YZDc-fmcmS-RCfa3e { transition: left 0.218s ease-out 0s, top 0.218s ease-out 0s, height 0.218s ease-out 0s, width 0.218s ease-out 0s; }

.ndfHFb-c4YZDc-fmcmS, .ndfHFb-c4YZDc-fmcmS-s2gQvd { bottom: 0px; position: absolute; top: 0px; width: 100%; }

.ndfHFb-c4YZDc-fmcmS-haAclf { height: 100%; position: absolute; width: 100%; }

.ndfHFb-c4YZDc-fmcmS-s2gQvd { overflow: auto; }

.ndfHFb-c4YZDc-fmcmS-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd { right: initial; }

.ndfHFb-c4YZDc-fmcmS-b0t70b { position: absolute; }

.ndfHFb-c4YZDc-fmcmS-bN97Pc { user-select: text; border: 20px solid transparent; font-family: "Courier New", Courier, monospace, arial, sans-serif; font-size: 14px; overflow-wrap: break-word; box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; background-color: rgb(255, 255, 255) !important; color: rgb(0, 0, 0) !important; }

.ndfHFb-c4YZDc-fmcmS-DARUcf { user-select: text; display: block; font-family: "Courier New", Courier, monospace, arial, sans-serif; margin: 0px; white-space: pre-wrap; overflow-wrap: break-word; background-color: rgb(255, 255, 255) !important; color: rgb(0, 0, 0) !important; }

.ndfHFb-c4YZDc-fmcmS-bN97Pc.ndfHFb-c4YZDc-fmcmS-kY93ue, .ndfHFb-c4YZDc-fmcmS-kY93ue .ndfHFb-c4YZDc-fmcmS-DARUcf { user-select: none; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf { height: 100%; position: absolute; width: 100%; z-index: 1; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q { position: absolute; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c { opacity: 0.2; background-color: rgb(34, 136, 255); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf { opacity: 0.5; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c { opacity: 0.4; background-color: rgb(52, 168, 83); }

.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-auswjd.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c { opacity: 1; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf:not([onclick]):not(:link):not(:visited) { background-color: transparent !important; }

.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf { opacity: 0.5; }

.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c { opacity: 0.4; background-color: rgb(251, 188, 4); }

.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-auswjd.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c { opacity: 1; }

.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b { display: none; }

.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-NowJzb { border-bottom: 2px solid rgb(251, 188, 4); }

.ndfHFb-c4YZDc-JUCs7e { border: 3px solid transparent; border-radius: 3px; display: inline-block; height: 63px; margin: 3px 0px 3px 3px; outline: none; width: 84px; }

.ndfHFb-c4YZDc-JUCs7e-SmKAyb { display: table-cell; height: inherit; vertical-align: middle; width: inherit; }

.ndfHFb-c4YZDc-JUCs7e img { display: block; margin: auto; }

.ndfHFb-c4YZDc-JUCs7e-Bz112c { width: 63px; height: 63px; }

.ndfHFb-c4YZDc-JUCs7e-RJLb9c { max-height: 63px; max-width: 84px; }

.ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-gk6SMd { border-color: transparent; }

.ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-ZmdkE, .ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-XpnDCe { border-color: rgb(156, 156, 156); }

.ndfHFb-c4YZDc-q77wGc { position: absolute; left: 50%; margin-right: -50%; transform: translate(-50%); border-radius: 3px; bottom: 12px; z-index: 3; overflow: hidden; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-q77wGc { border-radius: 100px; display: flex; }

.ndfHFb-c4YZDc-q77wGc .ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb, .ndfHFb-c4YZDc-q77wGc .ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb { background: rgba(0, 0, 0, 0.75); }

.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-C7uZwb-ibnC6b-Btuy5e { border-radius: 25%; padding: 0px; }

.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b .ndfHFb-c4YZDc-C7uZwb-ibnC6b-Btuy5e .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c { transform: scale(0.66667) translateY(-2px); }

.ndfHFb-c4YZDc-GSQQnc-LgbsSe, .ndfHFb-c4YZDc-MZArnb-LgbsSe, .ndfHFb-c4YZDc-TvD9Pc-LgbsSe { z-index: 1; min-height: 24px; }

.ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { opacity: 0.87; position: relative; margin-left: auto; margin-right: auto; }

.ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-GSQQnc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-MZArnb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c, .ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { height: 21px; width: 21px; margin-top: 3px; }

.ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px 0px; }

.ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1160px; }

.ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1280px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1528px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -1712px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c { background-position: 0px -2304px; height: 24px; width: 24px; margin: 0px; }

.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b .ndfHFb-c4YZDc-GSQQnc-LgbsSe { margin-left: 0px; }

.ndfHFb-c4YZDc-tk3N6e-suEOdc.tk3N6e-suEOdc { background-color: rgb(0, 0, 0); border-color: rgb(0, 0, 0); font-family: arial, sans-serif; z-index: 210; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tk3N6e-suEOdc.tk3N6e-suEOdc { border-radius: 2px; font-family: "Google Sans", Roboto, arial, sans-serif; }

.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-color: rgb(0, 0, 0) transparent; }

.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG, .ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG { border-color: transparent rgb(0, 0, 0); }

.ndfHFb-c4YZDc-neVct-RCfa3e { transition-property: left, top, width, height; transition-duration: 0.218s; transition-timing-function: cubic-bezier(0, 0, 0.2, 1); }

.ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e { transition-property: left, right, top, bottom; transition-duration: 0.218s; transition-timing-function: cubic-bezier(0, 0, 0.2, 1); }

.ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b { display: inline-block; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b { border: 1px solid transparent; border-radius: 2px; background: rgba(0, 0, 0, 0.75); margin: 0px; white-space: nowrap; }

.ndfHFb-c4YZDc-zM6fo-GMvhG-Bz112c { background-position: 0px -2584px; height: 18px; width: 18px; margin: 2px 4px; position: absolute; }

.ndfHFb-c4YZDc-zM6fo-GMvhG-fmcmS { line-height: 22px; margin: 2px 15px 2px 24px; font-size: 14px; font-weight: normal; }

.ndfHFb-c4YZDc-aTv5jf { border: 10px solid transparent; position: absolute; z-index: 0; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf { border: none; }

.ndfHFb-c4YZDc-aTv5jf-uquGtd { position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; z-index: 1; }

.ndfHFb-c4YZDc-aTv5jf-AHe6Kc { position: absolute; width: 100%; height: 100%; top: 0px; left: 0px; z-index: 1; }

.ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf { font: 13px arial; text-align: center; z-index: 2; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf a { text-decoration: underline; color: rgb(255, 255, 255) !important; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf { color: rgb(30, 30, 30); }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf a { color: rgb(30, 30, 30) !important; }

.ndfHFb-c4YZDc-aTv5jf-bVEB4e { background-color: black; cursor: pointer; position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; z-index: 2; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf-NziyQe-Bz112c:not(:link):not(:visited) { background-repeat: no-repeat; height: 77px; width: 77px; opacity: 0.8; background-image: url("//ssl.gstatic.com/s2/tt/images/play-overlay.png") !important; background-color: transparent !important; }

.ndfHFb-c4YZDc-aTv5jf-NziyQe-LgbsSe { z-index: 3; opacity: 0.8; position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc-aTv5jf-bVEB4e-RJLb9c { height: 100%; width: 100%; }

.ndfHFb-c4YZDc:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-aTv5jf-AHe6Kc { box-shadow: rgba(0, 0, 0, 0.35) 0px 4px 15px 2px; }

.ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde { position: absolute; top: 50%; left: 50%; margin-right: -50%; transform: translate(-50%, -50%); }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { background-image: url("//ssl.gstatic.com/docs/common/v-spinner_dark.gif") !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited) { background-image: none !important; }

.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS { color: rgb(255, 255, 255) !important; }

.ndfHFb-c4YZDc-LSZ0mb-fmcmS { margin-left: 5px; }

.ndfHFb-c4YZDc-LSZ0mb-hFsbo { border-left: 4px solid transparent; border-right: 4px solid transparent; margin-bottom: 1px; margin-left: 11px; display: inline-block; }

.ndfHFb-c4YZDc-LSZ0mb-hFsbo-hgHJW { border-top: 4px solid rgba(255, 255, 255, 0.87); }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-LSZ0mb-hFsbo-hgHJW { border-top: 4px solid rgb(255, 255, 255); }

.ndfHFb-c4YZDc-LSZ0mb-hFsbo-yHKmmc { border-bottom: 4px solid rgba(255, 255, 255, 0.87); }

.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-LSZ0mb-hFsbo-yHKmmc { border-bottom: 4px solid rgb(255, 255, 255); }

.ndfHFb-c4YZDc-kODWGd-xlL3N { height: 100%; position: absolute; left: auto; right: 10px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-LgbsSe { left: -35px; right: auto; position: absolute; top: 2px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c, .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c, .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c, .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c { height: 28px; width: 31px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c { background-position: 0px -2120px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c { background-position: 0px -2040px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c { background-position: 0px -560px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c { background-position: 0px -1400px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c { background-position: 0px -1408px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c { background-position: 0px -3794px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c { background-position: 0px -2810px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c { background-position: 0px -936px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-SxecR { width: 40px; }

.ndfHFb-c4YZDc-kODWGd-xlL3N-SxecR-PFprWc { height: 12px; width: 12px; }

.ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc { background: rgb(66, 133, 244); border-radius: 2px; color: rgb(0, 0, 0); font: 13px / 20px arial, sans-serif; position: absolute; width: 562px; z-index: 101; }

.ndfHFb-c4YZDc-deA65-di8rgd-LgbsSe { background: transparent; border: none; color: white; cursor: pointer; float: right; font-size: 14px; margin-bottom: auto; margin-left: auto; margin-top: auto; padding: 10px 16px; text-decoration: none; text-transform: uppercase; }

.ndfHFb-c4YZDc-deA65-di8rgd-LgbsSe:hover { outline: white auto 5px; }

.ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc-r4nke-fmcmS, .ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc-bN97Pc { float: left; font-size: 14px; font-weight: 500; padding: 10px 32px 10px 16px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb, .ndfHFb-c4YZDc-nJjxad-b0t70b { display: inline-block; white-space: nowrap; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb { height: 40px; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-b0t70b { margin-left: 10px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-Bz112c { opacity: 0.87; height: 21px; width: 21px; position: relative; margin-left: auto; margin-right: auto; margin-top: 3px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-Bz112c { opacity: 1; height: 24px; width: 24px; margin: 0px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-Bz112c { opacity: 0.47; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Bz112c { opacity: 1; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE { background-color: rgb(97, 97, 97); background-image: none; }

.ndfHFb-c4YZDc-nJjxad-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -2440px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -776px; }

.ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1360px; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1016px; }

.ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited) { background-position: 0px center; background-image: url("//ssl.gstatic.com/docs/common/v-spinner_dark.gif") !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited) { opacity: 1; background-image: none !important; }

.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-aZ2wEe { display: block; }

.ndfHFb-c4YZDc-nJjxad-SxecR { display: inline-block; height: 8px; margin-right: 10px; width: 100px; }

.ndfHFb-c4YZDc-nJjxad-SxecR .ndfHFb-c4YZDc-SxecR-skjTt-j4LONd { background-image: -webkit-linear-gradient(top, rgb(195, 195, 195), rgb(217, 217, 217)); background-color: rgb(217, 217, 217) !important; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-SxecR .ndfHFb-c4YZDc-SxecR-skjTt-j4LONd { background-image: none; box-shadow: rgba(0, 0, 0, 0.35) 0px 1px 1px 0px; background-color: rgb(255, 255, 255) !important; border-color: transparent !important; }

.ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc { background-image: -webkit-linear-gradient(top, rgb(0, 0, 0), rgb(48, 48, 48)); box-shadow: rgb(255, 255, 255) 0px 0px 5px 0px; border-radius: 6px; top: 18px; height: 10px; width: 10px; border: 1px solid rgb(255, 255, 255); background-color: rgb(21, 21, 21) !important; }

.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc { top: 16px; }

.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc { background-image: none; height: 8px; width: 8px; border: 2px solid rgb(255, 255, 255); margin-left: 10px; box-shadow: rgba(0, 0, 0, 0.35) 0px 1px 1px 0px; background-color: rgb(88, 89, 91) !important; }

.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-SxecR-PFprWc.ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc { background-image: none; box-shadow: rgba(30, 53, 69, 0.9) 0px 1px 1px 0px; background-color: rgb(255, 255, 255) !important; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb { display: inline-block; padding: 2px; vertical-align: middle; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { border-radius: 1px; width: 24px; height: 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe { border-radius: 100px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me { opacity: 0.47; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe .ndfHFb-c4YZDc-Bz112c { width: 24px; height: 24px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-m9bMae-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -2200px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-bEDTcc-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -552px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe .ndfHFb-c4YZDc-Bz112c { background-position: 0px -776px; }

.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe.ndfHFb-c4YZDc-nJjxad-S9gUrf .ndfHFb-c4YZDc-Bz112c { background-position: 0px -1016px; }

.EDlbXc-RTRLOc-OUyo8b { position: absolute; top: -1000px; height: 1px; overflow: hidden; }

.IyROMc-euCgFf-LJSvSb { background-image: url("//ssl.gstatic.com/docs/documents/share/images/sprite-24.svg"); }

.tk3N6e-cXJiPb { border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; transition: all 0s linear 1s, opacity 1s ease 0s; border-style: solid; border-width: 0px; font-size: 11px; height: 0px; opacity: 0; visibility: hidden; overflow: hidden; padding: 0px; text-align: center; }

.tk3N6e-cXJiPb-Tswv1b { background-color: rgb(249, 237, 190); border-color: rgb(240, 195, 109); color: rgb(51, 51, 51); }

.tk3N6e-cXJiPb-u0pjoe { background-color: rgb(72, 72, 72); border-color: rgb(32, 32, 32); color: rgb(255, 255, 255); }

.tk3N6e-cXJiPb-EfADOe { background-color: rgb(214, 233, 248); border-color: rgb(77, 144, 240); color: rgb(51, 51, 51); }

.tk3N6e-cXJiPb-GMvhG { background-color: rgb(221, 75, 57); border-color: rgb(96, 32, 25); color: rgb(255, 255, 255); }

.tk3N6e-cXJiPb-TSZdd { transition: opacity 0.218s ease 0s; border-width: 1px; min-height: 14px; height: auto; opacity: 1; visibility: visible; padding: 6px 16px; }

.tk3N6e-cXJiPb-yolsp.tk3N6e-cXJiPb-TSZdd { padding: 2px 16px; }

.euCgFf-X3SwIb-haAclf { font-family: Roboto, arial, sans-serif; font-size: 13px; font-weight: bold; position: fixed; display: inline-block; padding-bottom: 5px; }

.euCgFf-CJXtmf-Sx9Kwc .euCgFf-X3SwIb-haAclf { font-family: arial, sans-serif; }

.euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd { height: 21px; }

.euCgFf-X3SwIb-ma6Yeb { top: 23px; }

.euCgFf-X3SwIb-L7wHw { z-index: 3021; }

.euCgFf-PLEiK-Bz112c { opacity: 0.55; display: inline-block; width: 21px; height: 21px; margin-bottom: 1px; margin-top: 1px; margin-right: 1px; vertical-align: middle; }

.euCgFf-PLEiK-Ne3sFf, .euCgFf-PLEiK-hSRGPd { line-height: 21px; }

.euCgFf-PLEiK-hSRGPd, .euCgFf-PLEiK-hSRGPd:visited { color: rgb(17, 85, 204); text-decoration: none; cursor: pointer; }

.euCgFf-PLEiK-hSRGPd:focus { outline: none; }

.euCgFf-PLEiK-hSRGPd:active { color: rgb(209, 72, 54); }

.euCgFf-PLEiK-hSRGPd:disabled { color: rgb(34, 34, 34); cursor: default; }

.euCgFf-PLEiK-jCCvxc-Bz112c { background-position: 0px -212px; }

.euCgFf-PLEiK-Q8isyc-GEUYHe-Bz112c { background-position: 0px -778px; }

.euCgFf-PLEiK-iyXyEd-hSRGPd-Bz112c { background-position: 0px -412px; }

.VIpgJd-xl07Ob { border-radius: 0px; box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; transition: opacity 0.218s ease 0s; background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.2); cursor: default; font-size: 13px; margin: 0px; outline: none; padding: 6px 0px; position: absolute; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-linear-gradient(top, rgb(245, 245, 245), rgb(241, 241, 241)); border: 1px solid rgb(220, 220, 220); color: rgb(68, 68, 68); cursor: default; font-size: 11px; font-weight: bold; line-height: 27px; list-style: none; margin: 0px 2px; min-width: 46px; outline: none; padding: 0px 18px 0px 6px; text-align: center; text-decoration: none; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { background-color: rgb(255, 255, 255); border-color: rgb(243, 243, 243); color: rgb(184, 184, 184); }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; border-color: rgb(198, 198, 198); color: rgb(51, 51, 51); }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { border-color: rgb(77, 144, 254); }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-linear-gradient(top, rgb(238, 238, 238), rgb(224, 224, 224)); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); z-index: 2; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { vertical-align: top; white-space: nowrap; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(119, 119, 119) transparent; border-style: solid; border-width: 4px 4px 0px; height: 0px; width: 0px; position: absolute; right: 5px; top: 12px; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c { margin-top: -3px; opacity: 0.55; vertical-align: middle; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-gk6SMd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c { opacity: 0.9; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-gk6SMd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(89, 89, 89) transparent; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-qwU8Me { z-index: 1; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { z-index: 0; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-qwU8Me:focus, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-qwU8Me { z-index: 2; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu:focus, .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-LK5yu { z-index: 2; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-LK5yu { margin-left: -1px; border-bottom-left-radius: 0px; border-top-left-radius: 0px; min-width: 0px; padding-left: 0px; vertical-align: top; }

.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-qwU8Me { margin-right: 0px; border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.VIpgJd-j7LFlb, .VIpgJd-pWKtN, .VIpgJd-SFgmFf { position: relative; color: rgb(51, 51, 51); cursor: pointer; list-style: none; margin: 0px; padding: 6px 8em 6px 30px; white-space: nowrap; }

.VIpgJd-xl07Ob-RDtZlf .VIpgJd-j7LFlb, .VIpgJd-xl07Ob-GP8zAc .VIpgJd-j7LFlb { padding-left: 16px; vertical-align: middle; }

.VIpgJd-xl07Ob-KEZkZ .VIpgJd-j7LFlb { padding-right: 44px; }

.VIpgJd-j7LFlb-OWB6Me { cursor: default; }

.VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-x29Bmf, .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-bN97Pc { color: rgb(204, 204, 204) !important; }

.VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-Bz112c { opacity: 0.3; }

.VIpgJd-j7LFlb-sn54Q, .VIpgJd-j7LFlb-ZmdkE { background-color: rgb(238, 238, 238); border-color: rgb(238, 238, 238); border-style: dotted; border-width: 1px 0px; padding-top: 5px; padding-bottom: 5px; }

.VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-bN97Pc, .VIpgJd-j7LFlb-ZmdkE .VIpgJd-j7LFlb-bN97Pc { color: rgb(51, 51, 51); }

.VIpgJd-j7LFlb-MPu53c, .VIpgJd-j7LFlb-Bz112c { background-repeat: no-repeat; height: 21px; left: 3px; position: absolute; right: auto; top: 3px; vertical-align: middle; width: 21px; }

.VIpgJd-wQNmvb-gk6SMd { background-image: url("//ssl.gstatic.com/ui/v1/menu/checkmark.png"); background-repeat: no-repeat; background-position: left center; }

.VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-bN97Pc { color: rgb(51, 51, 51); }

.VIpgJd-j7LFlb-x29Bmf { color: rgb(119, 119, 119); direction: ltr; left: auto; padding: 0px 6px; position: absolute; right: 0px; text-align: right; }

.VIpgJd-j7LFlb-PQTlnb-brjg8b { text-decoration: underline; }

.VIpgJd-j7LFlb-PQTlnb-hgDUwe { color: rgb(119, 119, 119); font-size: 12px; padding-left: 4px; }

.VIpgJd-gqMrKb { border-top: 1px solid rgb(235, 235, 235); margin-top: 6px; margin-bottom: 6px; }

.euCgFf-CJXtmf-Sx9Kwc { overflow: auto; box-sizing: border-box; max-height: 100% !important; width: auto !important; }

* html .euCgFf-CJXtmf-Sx9Kwc { max-height: none !important; overflow: visible !important; }

:first-child + html .euCgFf-CJXtmf-Sx9Kwc { max-height: none !important; overflow: visible !important; }

.euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc, .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { padding: 0px; }

.euCgFf-CJXtmf-Sx9Kwc .euCgFf-CJXtmf-Sx9Kwc-L6cTce-r4nke { height: 0px; margin: 0px; padding: 0px; }

.euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { font-family: arial, sans-serif; font-weight: normal; }

.euCgFf-CJXtmf-bN97Pc-L5Fo6c { display: flex; height: 100%; width: 100%; border: none; }

.euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd { display: none; }

.euCgFf-CJXtmf-u0pjoe-Sx9Kwc { font-family: arial, sans-serif; font-size: 12px; width: 400px; z-index: 3000; }

.euCgFf-CJXtmf-ge6pde-BPrWId { height: 99px; text-align: center; width: 454px; }

.euCgFf-CJXtmf-aZ2wEe { background-image: url("//ssl.gstatic.com/docs/documents/share/images/spinner-1.gif"); display: inline-block; margin-top: 41px; width: 16px; height: 16px; }

.TzA9Ye-euCgFf-vWsuo-jOfkMb { font-size: 12pt; font-weight: bold; height: 19px; padding: 5px 10px; background-color: rgb(241, 244, 255); }

.TzA9Ye-euCgFf-vWsuo-bF1uUb { position: absolute; z-index: 150; background-color: rgb(255, 255, 255); opacity: 0; }

.euCgFf-CJXtmf-b0t70b-Sx9Kwc-euCgFf { height: 100%; width: 100%; }

.euCgFf-CJXtmf-b0t70b-Sx9Kwc-bF1uUb { position: absolute; z-index: 150; }

.euCgFf-CJXtmf-ynRLnc { position: absolute !important; left: -10000px !important; top: -10000px !important; }

.euCgFf-CJXtmf-ge6pde-Sx9Kwc { font-family: arial, sans-serif; z-index: 3000; }

.euCgFf-CJXtmf-E90Ek { display: none; position: absolute; bottom: 0px; right: 0px; color: rgb(119, 119, 119); font-size: 10px; }

.J2xVie-ndfHFb-euCgFf-CJXtmf-Sx9Kwc { border: none; border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.14) 0px 24px 38px 3px, rgba(0, 0, 0, 0.12) 0px 9px 46px 8px, rgba(0, 0, 0, 0.2) 0px 11px 15px -7px; padding: 0px; }

.Vkfede-uMX1Ee-euCgFf-CJXtmf-Sx9Kwc { height: 100vh; overflow: hidden; background-color: transparent !important; border: none !important; padding: 0px !important; width: 100vw !important; }

.Vkfede-uMX1Ee-euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { background: transparent; height: 100%; width: 100%; }

.XKSfm-Sx9Kwc.euCgFf-CJXtmf-Sx9Kwc.J2xVie-ndfHFb-euCgFf-CJXtmf-Sx9Kwc { padding: 0px; }

.Vkfede-uMX1Ee-euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke, .J2xVie-ndfHFb-euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { display: none; }

.tk3N6e-suEOdc { z-index: 30000; }

.zAYgkb-haAclf, .zAYgkb-Bz112c { display: inline-block; }

.zAYgkb-LgbsSe-Bz112c { margin: -3px 2px 0px -5px; vertical-align: middle !important; }

.zAYgkb-suEOdc-BPrWId { color: rgb(255, 255, 255); font-size: 13px; max-width: 300px; }

.zAYgkb-suEOdc-r4nke { font-size: 14px; font-weight: bold; }

.zAYgkb-suEOdc-fmcmS { font-weight: normal; }

.zAYgkb-suEOdc-Bz112c-haAclf { width: 25px; vertical-align: top; }

.zAYgkb-suEOdc-hgDUwe { border-top: 1px solid rgb(85, 85, 85); margin: 2px 0px; }

.tk3N6e-LgbsSe-n2to0e .zAYgkb-LgbsSe-Bz112c { opacity: 0.55; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-barxie .zAYgkb-LgbsSe-Bz112c, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-gk6SMd .zAYgkb-LgbsSe-Bz112c, .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE .zAYgkb-LgbsSe-Bz112c { opacity: 0.9; }

.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me .zAYgkb-LgbsSe-Bz112c { opacity: 0.333; }

.zAYgkb-g30GS-Bz112c-HLvlvd, .zAYgkb-d1sa2c-Bz112c-HLvlvd, .zAYgkb-QIk5de-g30GS-Bz112c-HLvlvd, .zAYgkb-QIk5de-d1sa2c-Bz112c-HLvlvd, .zAYgkb-BiKSr-PoC6nf-Bz112c-HLvlvd, .zAYgkb-IsSuNc-Bz112c-HLvlvd, .zAYgkb-UJflGc-Bz112c-HLvlvd, .zAYgkb-jsmBPd-Bz112c { width: 21px; height: 21px; background-repeat: no-repeat; vertical-align: bottom; }

.zAYgkb-g30GS-Oq668, .zAYgkb-pGuBYc-Oq668, .zAYgkb-QIk5de-Oq668, .zAYgkb-GEUYHe-Oq668, .zAYgkb-GMvhG-Oq668, .zAYgkb-iyXyEd-htvI8d-Oq668 { height: 18px; width: 18px; }

.zAYgkb-g30GS-Bz112c-HLvlvd { background-position: 0px -45px; }

.zAYgkb-d1sa2c-Bz112c-HLvlvd { background-position: 0px -562px; }

.zAYgkb-QIk5de-g30GS-Bz112c-HLvlvd { background-position: 0px -1004px; }

.zAYgkb-QIk5de-d1sa2c-Bz112c-HLvlvd { background-position: 0px -709px; }

.zAYgkb-BiKSr-PoC6nf-Bz112c-HLvlvd { background-position: 0px -932px; }

.zAYgkb-IsSuNc-Bz112c-HLvlvd { background-position: 0px -586px; }

.zAYgkb-UJflGc-Bz112c-HLvlvd { background-position: 0px -332px; }

.zAYgkb-jsmBPd-Bz112c { background-position: 0px -436px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-g30GS-Bz112c-HLvlvd { background-position: 0px -161px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-d1sa2c-Bz112c-HLvlvd { background-position: 0px -412px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-QIk5de-g30GS-Bz112c-HLvlvd { background-position: 0px -980px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-QIk5de-d1sa2c-Bz112c-HLvlvd { background-position: 0px -610px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-BiKSr-PoC6nf-Bz112c-HLvlvd { background-position: 0px -778px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-IsSuNc-Bz112c-HLvlvd { background-position: 0px 0px; }

.HB1eCd-n7vHCb-arrpzb .zAYgkb-UJflGc-Bz112c-HLvlvd { background-position: 0px -634px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-g30GS-Oq668 { background-position: 0px -236px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-pGuBYc-Oq668 { background-position: 0px -69px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-QIk5de-Oq668 { background-position: 0px -757px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-GEUYHe-Oq668 { background-position: 0px -24px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-GMvhG-Oq668 { background-position: 0px -90px; }

.HB1eCd-MqDS2b-uoC0bf .zAYgkb-suEOdc-r4nke, .HB1eCd-MqDS2b-uoC0bf .zAYgkb-suEOdc-fmcmS { color: rgb(242, 242, 242); font-size: 12px; font-weight: 400; }

.zAYgkb-iyXyEd-htvI8d-Oq668 { background-position: 0px -909px; }

.auswjd-mzNpsf-Sx9Kwc { background: rgb(255, 255, 255); border: 1px solid transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; position: absolute; z-index: 1003; padding: 24px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { font-size: 16px; position: relative; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-fmcmS { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 22px; font-weight: 400; line-height: 28px; display: inline-block; min-width: 200px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { color: rgb(60, 64, 67); }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; display: flex; justify-content: flex-end; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button { margin: 0px 0px 0px 12px; cursor: pointer; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button[disabled] { cursor: default; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button:first-child { margin-left: 0px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); border: 1px solid rgb(218, 220, 224) !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button:hover { background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button:focus { background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button:hover:focus { background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd button[disabled] { background: white; color: rgb(60, 64, 67); opacity: 0.38; border: 1px solid rgb(241, 243, 244) !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); border: 1px solid transparent !important; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover:focus { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active, .auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus:active { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; }

.auswjd-mzNpsf-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled] { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; }

.lZ2Ukb-Ujd07d-DARUcf-haAclf { left: 50%; margin: auto; position: absolute; top: 30%; transform: translate(-50%, -50%); width: 60%; }

.lZ2Ukb-Ujd07d-ndfHFb-r4nke-haAclf { align-items: center; display: inline-flex; margin: 0px 6px; }

.lZ2Ukb-Ujd07d-ndfHFb-r4nke { align-items: center; color: rgb(95, 99, 104); display: flex; font-family: "Google Sans"; font-size: 18px; font-style: normal; height: 16px; line-height: 23px; margin: 0px 6px; }

.lZ2Ukb-Ujd07d-ndfHFb-r4nke .lZ2Ukb-Ujd07d-ndfHFb-r4nke-jcJzye { font-weight: 500; margin-right: 3px; }

.lZ2Ukb-Ujd07d-Ne3sFf-haAclf { display: flex; height: 140px; margin-top: 60px; }

.lZ2Ukb-Ujd07d-r4nke { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1.75rem; font-weight: 400; letter-spacing: 0px; line-height: 2.25rem; color: rgb(32, 33, 36); margin-bottom: 8px; }

.lZ2Ukb-Ujd07d-nupQLb-Ne3sFf { font-style: normal; font-weight: normal; }

.lZ2Ukb-Ujd07d-ij8cu { color: rgb(95, 99, 104); font-family: Roboto; font-size: 14px; letter-spacing: 0.2px; line-height: 20px; }

.lZ2Ukb-Ujd07d-u0pjoe-xPjCTc { color: rgb(217, 48, 37); }

.lZ2Ukb-Ujd07d-Hn6s1b { margin-bottom: 20px; }

.lZ2Ukb-Bz112c { margin-right: 15px; }

.jcJzye-ndfHFb-Bz112c { background-repeat: no-repeat; height: 25px; width: 25px; }

.lZ2Ukb-E90Ek-Sx9Kwc-bN97Pc { max-height: 640px; max-width: 1024px; overflow: auto; }

.KCJqBf-Sx9Kwc-bN97Pc { max-height: 428px; max-width: 1024px; overflow: auto; }

.KCJqBf-O0r3Gd-Sx9Kwc { height: 512px; }

#apps-debug-tracers { display: none; }

.ndfHFb-c4YZDc-E90Ek-haAclf { margin-bottom: 6px; margin-right: 6px; vertical-align: top; }

.HB1eCd-E90Ek-Tswv1b, .HB1eCd-E90Ek-Tswv1b a { font-size: 8px; color: rgb(119, 119, 119) !important; }

.ndfHFb-c4YZDc-E90Ek-haAclf.HB1eCd-E90Ek-Tswv1b { display: flex; position: absolute; right: 0px; bottom: 0px; z-index: 300; }

.lZ2Ukb-zzT4b-PGTmtf { border-style: solid; border-width: 1px; font-size: 12px; margin-bottom: 14px; padding: 12px; }

.ndfHFb-c4YZDc-uoC0bf .lZ2Ukb-zzT4b-PGTmtf { background: rgb(255, 223, 153); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 14px; line-height: 20px; border-radius: 4px; }

.lZ2Ukb-zzT4b-ij8cu { color: rgb(90, 90, 90); font-size: 12px; height: 16px; margin-bottom: 5px; overflow: hidden; }

.ndfHFb-c4YZDc-uoC0bf .lZ2Ukb-zzT4b-ij8cu { height: 30px; font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 14px; line-height: 20px; color: rgb(227, 227, 227); }

.lZ2Ukb-zzT4b-B7I4Od { border-color: rgb(204, 204, 204); direction: ltr; font-size: 12px; height: 100%; margin-bottom: 5px; overflow: auto; resize: none; width: 100%; }

.ndfHFb-c4YZDc-uoC0bf .lZ2Ukb-zzT4b-B7I4Od { margin: 0px; width: auto; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc { background: rgb(31, 31, 31); padding: 24px; border-radius: 8px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { background-color: rgb(31, 31, 31); color: rgb(227, 227, 227); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 24px; line-height: 32px; margin: 0px 0px 24px; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc { display: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc { background-color: rgb(31, 31, 31); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 16px; line-height: 24px; display: flex; flex-direction: column; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc .XKSfm-Sx9Kwc-c6xFrd { margin: 24px 0px 0px 24px; border-radius: 100px; background: rgb(31, 31, 31); color: rgb(168, 199, 250); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 500; font-size: 14px; line-height: 20px; border: none; display: flex; justify-content: flex-end; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc button { margin: 0px 0px 0px 24px; border-radius: 100px; background: rgb(31, 31, 31); color: rgb(168, 199, 250); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 500; font-size: 14px; line-height: 20px; border: none; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc button:hover { background: rgba(168, 199, 250, 0.08); color: rgb(168, 199, 250); border: none; }

.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc button:focus, .ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-e1YmVc-Sx9Kwc button:active { background: rgba(168, 199, 250, 0.12); color: rgb(168, 199, 250); border: none; outline: none; box-shadow: none; }

body { font-family: Roboto, sans-serif; }

.XKSfm-Sx9Kwc { z-index: 102; }

.XKSfm-Sx9Kwc-xJ5Hnf { z-index: 101; }

.Chn84b-haAclf { left: 0px; top: 0px; background-color: transparent; border: none; height: 100%; width: 100%; overflow: hidden; padding: 0px; position: absolute; z-index: 2500; }

.Chn84b-haAclf.xTMeO { display: none; }

.Chn84b-L5Fo6c-haAclf { height: 100%; width: 100%; background: transparent; padding: 0px; position: absolute; z-index: 1; }

.ge6pde .Chn84b-L5Fo6c-haAclf { opacity: 0; }

.Chn84b-o1DAbe-aZ2wEe-Lb81de { transform: translate(-50%, -50%); left: 50%; position: absolute; top: 50%; z-index: 1; }

.Chn84b-o1DAbe-ge6pde-haAclf-Lb81de { position: absolute; inset: 0px; overflow: hidden; border: none; padding: 0px; display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; background-color: var(--dt-scrim,rgba(32,33,36,.6)); visibility: hidden; z-index: 2; }

.ge6pde .Chn84b-o1DAbe-ge6pde-haAclf-Lb81de { visibility: visible; }

.Chn84b-o1DAbe-ge6pde-Sx9Kwc-Lb81de { width: 616px; height: 516px; max-width: 616px; max-height: 516px; min-width: 512px; min-height: 272px; border-radius: 8px; background-color: white; padding: 0px; margin: 20px; overflow: hidden; position: relative; }

.Chn84b-o1DAbe-ge6pde-fmcmS-Lb81de { color: rgba(32, 33, 36, 0.87); font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-headline-small-spacing,0); font-size: 24px; left: 24px; position: absolute; top: 22px; line-height: 32px; }

.Chn84b-o1DAbe-ge6pde-TvD9Pc-LgbsSe { background: url("https://fonts.gstatic.com/s/i/short-term/release/googlesymbols/close/default/24px.svg"); border: 0px; cursor: pointer; height: 24px; opacity: 0.87; position: absolute; right: 24px; top: 22px; width: 24px; }

.Chn84b-o1DAbe-ge6pde-TvD9Pc-suEOdc { visibility: hidden; border-radius: 2px; border: 0px; background-color: rgb(32, 33, 36); color: rgb(255, 255, 255); position: absolute; z-index: 1; right: 24px; top: 48px; opacity: 1; overflow-x: hidden; padding: 5px 8px 6px; text-align: center; font-size: 12px; }

.Chn84b-o1DAbe-ge6pde-TvD9Pc:hover .Chn84b-o1DAbe-ge6pde-TvD9Pc-suEOdc { visibility: visible; }

.oErxNe-pSzOP { width: 36px; height: 36px; overflow: hidden; animation: 1568.63ms linear 0s infinite normal none running mspin-rotate; }

.oErxNe-pSzOP .oErxNe-WkJb5 { animation: 5332ms steps(4) 0s infinite normal none running mspin-revrot; }

.oErxNe-pSzOP .oErxNe-aZ2wEe { background-image: url("//ssl.gstatic.com/docs/picker/images/loading_spinner.svg"); background-size: 100%; width: 11664px; height: 36px; animation: 5332ms steps(324) 0s infinite normal none running mspin-medium-film; }

@-webkit-keyframes mspin-medium-film { 
  0% { transform: translateX(0px); }
  100% { transform: translateX(-11664px); }
}

@keyframes mspin-medium-film { 
  0% { transform: translateX(0px); }
  100% { transform: translateX(-11664px); }
}

@-webkit-keyframes mspin-rotate { 
  0% { transform: rotate(0deg); }
  100% { transform: rotate(360deg); }
}

@keyframes mspin-rotate { 
  0% { transform: rotate(0deg); }
  100% { transform: rotate(360deg); }
}

@-webkit-keyframes mspin-revrot { 
  0% { transform: rotate(0deg); }
  100% { transform: rotate(-360deg); }
}

@keyframes mspin-revrot { 
  0% { transform: rotate(0deg); }
  100% { transform: rotate(-360deg); }
}

@keyframes mspin-medium-film { 
  0% { transform: translateX(0px); }
  100% { transform: translateX(-11664px); }
}

.ndfHFb-w37qKe-ppgLk-V68bde { display: flex; vertical-align: middle; }

.ndfHFb-w37qKe-ppgLk-V68bde-sfGayb-SKd3Ne { margin: auto; }

.ndfHFb-w37qKe-V68bde { position: absolute; z-index: 1002; box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; background-color: rgb(241, 241, 241); border: 1px solid rgba(0, 0, 0, 0.2); color: rgb(110, 110, 110); font-size: 13px; font-weight: normal; text-align: left; white-space: nowrap; }

.ndfHFb-w37qKe-V68bde-i5vt6e-L6cTce :focus { outline: none; }

.ndfHFb-w37qKe-V68bde-bN97Pc { display: flex; padding: 10px; }

.ndfHFb-w37qKe-V68bde-Ne3sFf { overflow: hidden; text-overflow: ellipsis; -webkit-box-orient: vertical; -webkit-line-clamp: 6; display: -webkit-box; max-height: 90px; margin: auto; max-width: 160px; padding-right: 10px; word-break: break-word; }

.ndfHFb-w37qKe-LgbsSe { display: inline-block; margin: auto; }

.ndfHFb-w37qKe-V68bde-hSRGPd-SKd3Ne { color: rgb(17, 85, 204); cursor: pointer; padding: 0px 7px; }

.ndfHFb-w37qKe-V68bde-TvD9Pc-SKd3Ne { cursor: pointer; height: 15px; padding: 3px; vertical-align: middle; }

.ndfHFb-w37qKe-V68bde-hSRGPd-SKd3Ne.ndfHFb-w37qKe-LgbsSe-ZmdkE { text-decoration: underline; }

.ndfHFb-w37qKe-V68bde-hFsbo { position: absolute; width: 20px; }

.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe, .ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc { content: ""; display: block; height: 0px; position: absolute; width: 0px; }

.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe { border: 10px solid; }

.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc { border: 9px solid; }

.ndfHFb-w37qKe-V68bde-Ya1KTb { bottom: 0px; }

.ndfHFb-w37qKe-V68bde-d6mlqf { top: -10px; }

.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe, .ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe { border-color: rgba(0, 0, 0, 0.2) transparent; left: 0px; }

.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc, .ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc { border-color: rgb(241, 241, 241) transparent; left: 1px; }

.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe, .ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc { border-bottom-width: 0px; }

.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe { border-top-width: 0px; }

.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc { border-top-width: 0px; top: 2px; }

.ndfHFb-w37qKe-Sx9Kwc { box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; background-image: ; background-position-x: ; background-position-y: ; background-size: ; background-repeat-x: ; background-repeat-y: ; background-attachment: ; background-origin: ; background-color: ; background-clip: padding-box; color: var(--dt-on-surface,#3c4043); font-family: inherit; outline: 0px; padding: 24px; position: absolute; width: 560px; z-index: 2204; }

.ndfHFb-w37qKe-Sx9Kwc-xJ5Hnf { background: var(--dt-on-surface,#3c4043); left: 0px; position: absolute; top: 0px; z-index: 2203; }

div.ndfHFb-w37qKe-Sx9Kwc-xJ5Hnf { opacity: 0.5; }

.ndfHFb-w37qKe-Sx9Kwc-r4nke { background-color: var(--dt-background,#fff); color: var(--dt-on-surface,#3c4043); cursor: default; font-size: 20px; font-weight: normal; line-height: 24px; }

.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc { height: 11px; margin: 24px; opacity: 0.7; padding: 6px; position: absolute; right: 0px; top: 0px; width: 11px; }

.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc::after { background: url("//ssl.gstatic.com/ui/v1/dialog/close-x.png"); content: ""; height: 11px; position: absolute; width: 11px; }

.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.ndfHFb-w37qKe-Sx9Kwc-bN97Pc { background-color: var(--dt-background,#fff); font-size: 16px; line-height: 1.4em; padding-top: 24px; padding-bottom: 24px; overflow-wrap: break-word; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd { text-align: right; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe { border-radius: 2px; background-color: var(--dt-surface-variant,#f1f3f4); background-image: linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1); border: 1px solid rgba(0, 0, 0, 0.1); color: var(--dt-on-surface,#3c4043); cursor: default; font-family: inherit; font-size: 11px; font-weight: bold; height: 29px; line-height: 27px; margin: 0px 0px 0px 16px; min-width: 72px; outline: 0px; padding: 0px 8px; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: var(--dt-surface-variant,#f1f3f4); background-image: linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1); border: 1px solid rgb(198, 198, 198); color: var(--dt-on-surface,#3c4043); }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:active { background-color: var(--dt-surface-variant,#f1f3f4); background-image: linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1); border: 1px solid rgb(198, 198, 198); color: var(--dt-on-surface,#3c4043); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:focus { border: 1px solid var(--dt-primary,#1a73e8); }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe[disabled] { box-shadow: none; background-position-x: ; background-position-y: ; background-size: ; background-repeat-x: ; background-repeat-y: ; background-attachment: ; background-origin: ; background-clip: ; background-color: ; background-image: none; border: 1px solid rgba(0, 0, 0, 0.5); color: rgba(0, 0, 0, 0.26); }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc { background-color: var(--dt-primary,#1a73e8); background-image: linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8)); border: 1px solid var(--dt-primary,#1a73e8); color: var(--dt-background,#fff); }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover { background-color: var(--dt-primary,#1a73e8); background-image: linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8)); border: 1px solid var(--dt-primary,#1a73e8); color: var(--dt-background,#fff); }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active { background-color: var(--dt-primary,#1a73e8); background-image: linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8)); border: 1px solid var(--dt-primary,#1a73e8); color: var(--dt-background,#fff); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled] { box-shadow: none; background: var(--dt-primary,#1a73e8); color: var(--dt-background,#fff); opacity: 0.5; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-xl07Ob { box-shadow: none; margin-bottom: -24px; padding: 0px; position: relative; z-index: inherit; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb { color: var(--dt-on-surface,#3c4043); font-size: 13px; height: 16px; margin: 0px; opacity: 0.87; padding: 0px 0px 24px 16px; }

.ndfHFb-w37qKe-Sx9Kwc-tlSJBe-V1ur5d { font-weight: bold; }

.ndfHFb-w37qKe-Sx9Kwc-rymPhb-ibnC6b { display: block; overflow: hidden; text-overflow: ellipsis; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-sn54Q { border-left: 0px; background-color: inherit; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-bN97Pc { margin: 0px; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-bN97Pc, .ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-bN97Pc { color: inherit; }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-auswjd .VIpgJd-j7LFlb-MPu53c { background: rgb(235, 235, 235); }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-AHmuwe .VIpgJd-j7LFlb-MPu53c { border-color: var(--dt-primary,#1a73e8); }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd { background: rgba(255, 255, 255, 0); }

.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-MPu53c::after { border-radius: 50%; background: rgb(96, 96, 96); content: ""; display: block; }

.ndfHFb-aZ2wEe { height: 44px; overflow: hidden; position: relative; }

.ndfHFb-vyDMJf-aZ2wEe { height: 28px; left: 50%; margin-left: -14px; position: absolute; top: 8px; width: 28px; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd { animation: 1568ms linear 0s infinite normal none running container-rotate; }

@-webkit-keyframes container-rotate { 
  100% { transform: rotate(360deg); }
}

@keyframes container-rotate { 
  100% { transform: rotate(360deg); }
}

.aZ2wEe-pbTTYe { position: absolute; width: 100%; height: 100%; opacity: 0; }

.aZ2wEe-v3pZbf { border-color: rgb(66, 133, 244); }

.aZ2wEe-oq6NAc { border-color: rgb(219, 68, 55); }

.aZ2wEe-gS7Ybc { border-color: rgb(244, 180, 0); }

.aZ2wEe-nllRtd { border-color: rgb(15, 157, 88); }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-v3pZbf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running blue-fade-in-out; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-oq6NAc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running red-fade-in-out; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-gS7Ybc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running yellow-fade-in-out; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-nllRtd { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running green-fade-in-out; }

@-webkit-keyframes fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@keyframes fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@-webkit-keyframes blue-fade-in-out { 
  0% { opacity: 1; }
  25% { opacity: 1; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 1; }
  100% { opacity: 1; }
}

@keyframes blue-fade-in-out { 
  0% { opacity: 1; }
  25% { opacity: 1; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 1; }
  100% { opacity: 1; }
}

@-webkit-keyframes red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 1; }
  50% { opacity: 1; }
  51% { opacity: 0; }
}

@keyframes red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 1; }
  50% { opacity: 1; }
  51% { opacity: 0; }
}

@-webkit-keyframes yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 1; }
  75% { opacity: 1; }
  76% { opacity: 0; }
}

@keyframes yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 1; }
  75% { opacity: 1; }
  76% { opacity: 0; }
}

@-webkit-keyframes green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 1; }
  90% { opacity: 1; }
  100% { opacity: 0; }
}

@keyframes green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 1; }
  90% { opacity: 1; }
  100% { opacity: 0; }
}

.aZ2wEe-pehrl-TpMipd { position: absolute; box-sizing: border-box; top: 0px; left: 45%; width: 10%; height: 100%; overflow: hidden; border-color: inherit; }

.aZ2wEe-pehrl-TpMipd .aZ2wEe-LkdAo { width: 1000%; left: -450%; }

.aZ2wEe-LkdAo-e9ayKc { display: inline-block; position: relative; width: 50%; height: 100%; overflow: hidden; border-color: inherit; }

.aZ2wEe-LkdAo-e9ayKc .aZ2wEe-LkdAo { width: 200%; }

.aZ2wEe-LkdAo { box-sizing: border-box; height: 100%; border-width: 3px; border-style: solid; border-top-color: inherit; border-right-color: inherit; border-left-color: inherit; border-radius: 50%; animation: 0s ease 0s 1 normal none running none; border-bottom-color: transparent !important; }

.aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { transform: rotate(129deg); border-right-color: transparent !important; }

.aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { left: -100%; transform: rotate(-129deg); border-left-color: transparent !important; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running left-spin; }

.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running right-spin; }

@-webkit-keyframes left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@keyframes left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@-webkit-keyframes right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@keyframes right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

.aZ2wEe-hj4D6d { position: absolute; inset: 0px; }

.wvGCSb-VkLyEc-Sx9Kwc { font-size: 14px; white-space: normal; width: 472px; }

.wvGCSb-VkLyEc-Sx9Kwc .wvGCSb-VkLyEc-Sx9Kwc-VdSJob { width: 424px; }

.wvGCSb-VkLyEc-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-bN97Pc { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.wvGCSb { color: black; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; white-space: normal; }

.wvGCSb.HB1eCd-UMrnmb { font-size: 14px; }

.wvGCSb .tk3N6e-LgbsSe { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe { margin: 0px 8px 0px 0px; min-width: 24px; vertical-align: middle; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgba(0, 0, 0, 0.06); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe-auswjd { box-shadow: none; background-color: rgba(0, 0, 0, 0.12); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: white; color: rgb(26, 115, 232); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(218, 220, 224) !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(241, 243, 244) !important; }

@media (forced-colors: active) {
  .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-XpnDCe { outline: highlight solid 1px; outline-offset: -4px; }
}

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(193, 216, 251) !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(204, 224, 252) !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { background: rgb(225, 236, 254); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(187, 212, 251) !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; height: 24px; padding: 3px 12px 5px; border: 1px solid transparent !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid transparent !important; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb .XKSfm-Sx9Kwc-r4nke { font-size: 16px; }

.HB1eCd-UMrnmb .wvGCSb .XKSfm-Sx9Kwc-r4nke { font-size: 22px; }

.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: normal; }

.HB1eCd-UMrnmb .lI7fHe-XKSfm.XKSfm-Sx9Kwc { width: 300px; }

.HB1eCd-UMrnmb .lI7fHe-XKSfm .XKSfm-Sx9Kwc-r4nke-fmcmS { display: block; width: 220px; overflow-wrap: break-word; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e, .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(11, 87, 208); color: white; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { background: white; color: rgb(11, 87, 208); border-color: rgb(199, 199, 199) !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { height: 36px; line-height: 16px; padding: 9px 16px; color: rgb(31, 31, 31); cursor: default; background: rgba(31, 31, 31, 0.12); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { height: 36px; line-height: 16px; padding: 9px 16px; background-color: rgba(11, 87, 208, 0.08); box-shadow: none; color: rgb(11, 87, 208); border-color: rgb(199, 199, 199) !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-auswjd { border-width: 1px; border-style: solid; border-image: initial; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background-color: rgba(11, 87, 208, 0.12); box-shadow: none; color: rgb(11, 87, 208); border-color: rgb(11, 87, 208) !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(228, 228, 228); color: rgb(31, 31, 31); cursor: default; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(41, 107, 214); color: white; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { height: 36px; line-height: 16px; padding: 9px 16px; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 2px 6px 2px; background: rgb(30, 100, 212); color: white; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe { background: none; border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-auswjd { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.HB1eCd-uoC0bf-fmcmS-LgbsSe { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; white-space: nowrap; color: rgb(11, 87, 208); padding: 9px 12px; }

.HB1eCd-uoC0bf-fmcmS-LgbsSe.HB1eCd-uoC0bf-LgbsSe-ZmdkE { color: rgb(11, 87, 208); padding: 9px 12px; background-color: rgba(11, 87, 208, 0.08); }

.HB1eCd-uoC0bf-fmcmS-LgbsSe.HB1eCd-uoC0bf-LgbsSe-XpnDCe { color: rgb(11, 87, 208); padding: 9px 12px; background-color: rgba(11, 87, 208, 0.12); outline: none; }

.HB1eCd-uoC0bf-fmcmS-LgbsSe.HB1eCd-uoC0bf-LgbsSe-OWB6Me { padding: 9px 12px; color: rgb(31, 31, 31); cursor: default; }

.HB1eCd-uoC0bf-MFS4be-LgbsSe { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; background: rgb(11, 87, 208); color: rgb(255, 255, 255); }

.HB1eCd-uoC0bf-MFS4be-LgbsSe.HB1eCd-uoC0bf-LgbsSe-ZmdkE { color: rgb(255, 255, 255); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 1px 3px 1px; background: rgb(31, 100, 212); }

.HB1eCd-uoC0bf-MFS4be-LgbsSe.HB1eCd-uoC0bf-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(40, 107, 214); outline: none; }

.HB1eCd-uoC0bf-MFS4be-LgbsSe.HB1eCd-uoC0bf-LgbsSe-auswjd { color: rgb(255, 255, 255); background: rgb(40, 107, 214); outline: none; }

.HB1eCd-uoC0bf-MFS4be-LgbsSe.HB1eCd-uoC0bf-LgbsSe-OWB6Me { background: rgba(31, 31, 31, 0.12); color: rgba(31, 31, 31, 0.38); cursor: default; }

.HB1eCd-uoC0bf-INsAgc-LgbsSe { border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; height: 40px; line-height: 20px; padding: 9px 24px; white-space: nowrap; border: 1px solid rgb(116, 119, 117); color: rgb(11, 87, 208); }

.HB1eCd-uoC0bf-INsAgc-LgbsSe.HB1eCd-uoC0bf-LgbsSe-ZmdkE { border: 1px solid rgb(116, 119, 117); color: rgb(11, 87, 208); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 1px 3px 1px; background: rgba(11, 87, 208, 0.08); }

.HB1eCd-uoC0bf-INsAgc-LgbsSe.HB1eCd-uoC0bf-LgbsSe-XpnDCe { color: rgb(11, 87, 208); background: rgba(11, 87, 208, 0.12); border: 1px solid rgb(11, 87, 208); outline: none; }

.HB1eCd-uoC0bf-INsAgc-LgbsSe.HB1eCd-uoC0bf-LgbsSe-auswjd { border: 1px solid rgb(116, 119, 117); color: rgb(11, 87, 208); background: rgba(11, 87, 208, 0.12); outline: none; }

.HB1eCd-uoC0bf-INsAgc-LgbsSe.HB1eCd-uoC0bf-LgbsSe-OWB6Me { border: 1px solid rgba(31, 31, 31, 0.12); color: rgba(31, 31, 31, 0.38); cursor: default; }

.HB1eCd-uoC0bf-LgbsSe { margin: 0px 4px; }

@media screen and (forced-colors: active) {
  .HB1eCd-uoC0bf-LgbsSe.HB1eCd-uoC0bf-LgbsSe-XpnDCe { outline: highlight solid 1px; outline-offset: -4px; }
}

.LgbsSe-bN97Pc-SfQLQb-fuEl3d-Q3DXx-Q4BLdf { display: flex; gap: 8px; }

.HB1eCd-HzV7m .LgbsSe-bN97Pc-SfQLQb-fuEl3d-Q3DXx-Q4BLdf .HB1eCd-Bz112c { margin: 0px; }

.LgbsSe-bN97Pc-pUia2e-SfQLQb-Bz112c { margin-left: -8px; }

.LgbsSe-bN97Pc-emzOGe-SfQLQb-Bz112c { margin-right: -8px; }

.HB1eCd-UMrnmb .HB1eCd-HzV7m .LgbsSe-bN97Pc-Bz112c-OWB6Me .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_dark.svg"); opacity: 0.38; }

.HB1eCd-Guievd-WqyaDf .HB1eCd-uoC0bf-MFS4be-LgbsSe .LgbsSe-bN97Pc-Bz112c-qnnXGd .HB1eCd-Bz112c-RJLb9c { filter: unset; }

.HB1eCd-uoC0bf-LgbsSe:not(.HB1eCd-uoC0bf-LgbsSe-OWB6Me) .LgbsSe-bN97Pc-Bz112c-OWB6Me, .HB1eCd-uoC0bf-LgbsSe-OWB6Me .LgbsSe-bN97Pc-Bz112c-qnnXGd { display: none; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc { background: rgb(255, 255, 255); border: 1px solid transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; position: absolute; z-index: 1003; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); left: 0px; position: absolute; top: 0px; z-index: 998; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc:focus { outline: none; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke { border-bottom: none; padding: 24px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-fmcmS { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 22px; font-weight: 400; line-height: 28px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { height: 24px; position: absolute; right: 24px; top: 26px; width: 24px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-bN97Pc { min-width: 312px; padding: 0px 24px 24px; color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-c6xFrd { display: flex; justify-content: flex-end; padding: 24px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe, .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe { text-transform: none; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-F75qrd-wcotoc-JIbuQc-LgbsSe.HB1eCd-HzV7m-LgbsSe { margin-left: 12px; }

.VfPpkd-JGcpL-uI4vCe-LkdAo, .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: var(--mdc-theme-primary,#6200ee); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .VfPpkd-JGcpL-uI4vCe-LkdAo, .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.VfPpkd-JGcpL-uI4vCe-u014N { stroke: transparent; }

@-webkit-keyframes mdc-circular-progress-container-rotate { 
  100% { transform: rotate(1turn); }
}

@keyframes mdc-circular-progress-container-rotate { 
  100% { transform: rotate(1turn); }
}

@-webkit-keyframes mdc-circular-progress-spinner-layer-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@keyframes mdc-circular-progress-spinner-layer-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@-webkit-keyframes mdc-circular-progress-color-1-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@keyframes mdc-circular-progress-color-1-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@-webkit-keyframes mdc-circular-progress-color-2-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
  100% { opacity: 0; }
}

@keyframes mdc-circular-progress-color-2-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
  100% { opacity: 0; }
}

@-webkit-keyframes mdc-circular-progress-color-3-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
  100% { opacity: 0; }
}

@keyframes mdc-circular-progress-color-3-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
  100% { opacity: 0; }
}

@-webkit-keyframes mdc-circular-progress-color-4-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes mdc-circular-progress-color-4-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@-webkit-keyframes mdc-circular-progress-left-spin { 
  0% { transform: rotate(265deg); }
  50% { transform: rotate(130deg); }
  100% { transform: rotate(265deg); }
}

@keyframes mdc-circular-progress-left-spin { 
  0% { transform: rotate(265deg); }
  50% { transform: rotate(130deg); }
  100% { transform: rotate(265deg); }
}

@-webkit-keyframes mdc-circular-progress-right-spin { 
  0% { transform: rotate(-265deg); }
  50% { transform: rotate(-130deg); }
  100% { transform: rotate(-265deg); }
}

@keyframes mdc-circular-progress-right-spin { 
  0% { transform: rotate(-265deg); }
  50% { transform: rotate(-130deg); }
  100% { transform: rotate(-265deg); }
}

.VfPpkd-JGcpL-P1ekSe { display: inline-flex; position: relative; direction: ltr; line-height: 0; transition: opacity 0.25s cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-JGcpL-uI4vCe-haAclf, .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G, .VfPpkd-JGcpL-IdXvz-haAclf, .VfPpkd-JGcpL-QYI5B-pbTTYe { position: absolute; width: 100%; height: 100%; }

.VfPpkd-JGcpL-uI4vCe-haAclf { transform: rotate(-90deg); }

.VfPpkd-JGcpL-IdXvz-haAclf { font-size: 0px; letter-spacing: 0px; white-space: nowrap; opacity: 0; }

.VfPpkd-JGcpL-uI4vCe-LkdAo-Bd00G, .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { fill: transparent; }

.VfPpkd-JGcpL-uI4vCe-LkdAo { transition: stroke-dashoffset 0.5s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-JGcpL-OcUoKf-TpMipd { position: absolute; top: 0px; left: 47.5%; box-sizing: border-box; width: 5%; height: 100%; overflow: hidden; }

.VfPpkd-JGcpL-OcUoKf-TpMipd .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { left: -900%; width: 2000%; transform: rotate(180deg); }

.VfPpkd-JGcpL-lLvYUc-e9ayKc { display: inline-flex; position: relative; width: 50%; height: 100%; overflow: hidden; }

.VfPpkd-JGcpL-lLvYUc-e9ayKc .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { width: 200%; }

.VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { left: -100%; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-uI4vCe-haAclf { opacity: 0; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf { opacity: 1; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf { animation: 1.56824s linear 0s infinite normal none running mdc-circular-progress-container-rotate; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-QYI5B-pbTTYe { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-spinner-layer-rotate; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-R6PoUb { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-spinner-layer-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-color-1-fade-in-out; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-ibL1re { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-spinner-layer-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-color-2-fade-in-out; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-c5RTEf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-spinner-layer-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-color-3-fade-in-out; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-II5mzb { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-spinner-layer-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-color-4-fade-in-out; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-LK5yu .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-left-spin; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running mdc-circular-progress-right-spin; }

.VfPpkd-JGcpL-P1ekSe-OWXEXe-xTMeO { opacity: 0; }

.VfPpkd-z59Tgd { border-radius: var(--mdc-shape-small,4px); }

.VfPpkd-Djsh7e-XxIAqe-ma6Yeb, .VfPpkd-Djsh7e-XxIAqe-cGMI2b { border-radius: var(--mdc-shape-small,4px); }

.VfPpkd-z59Tgd { color: var(--mdc-theme-text-primary-on-dark,white); }

.VfPpkd-z59Tgd { background-color: rgba(0, 0, 0, 0.6); }

.VfPpkd-MlC99b { color: var(--mdc-theme-text-primary-on-light,rgba(0,0,0,.87)); }

.VfPpkd-IqDDtd { color: rgba(0, 0, 0, 0.6); }

.VfPpkd-IqDDtd-hSRGPd { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd, .VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb, .VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b { background-color: rgb(255, 255, 255); }

.VfPpkd-z59Tgd { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-caption-font-size,.75rem); font-weight: var(--mdc-typography-caption-font-weight,400); letter-spacing: var(--mdc-typography-caption-letter-spacing,.0333333333em); text-decoration: var(--mdc-typography-caption-text-decoration,inherit); text-transform: var(--mdc-typography-caption-text-transform,inherit); }

.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 1px -2px, rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 1px 5px 0px; border-radius: 4px; line-height: 20px; }

.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-BFbNVe-bF1uUb { width: 100%; height: 100%; top: 0px; left: 0px; }

.VfPpkd-z59Tgd .VfPpkd-MlC99b { display: block; margin-top: 0px; -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle2-font-size,.875rem); line-height: var(--mdc-typography-subtitle2-line-height,1.375rem); font-weight: var(--mdc-typography-subtitle2-font-weight,500); letter-spacing: var(--mdc-typography-subtitle2-letter-spacing,.0071428571em); text-decoration: var(--mdc-typography-subtitle2-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle2-text-transform,inherit); }

.VfPpkd-z59Tgd .VfPpkd-MlC99b::before { display: inline-block; width: 0px; height: 24px; content: ""; vertical-align: 0px; }

.VfPpkd-z59Tgd .VfPpkd-IqDDtd { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-body2-font-size,.875rem); line-height: var(--mdc-typography-body2-line-height,1.25rem); font-weight: var(--mdc-typography-body2-font-weight,400); letter-spacing: var(--mdc-typography-body2-letter-spacing,.0178571429em); text-decoration: var(--mdc-typography-body2-text-decoration,inherit); text-transform: var(--mdc-typography-body2-text-transform,inherit); }

.VfPpkd-z59Tgd { word-break: var(--mdc-tooltip-word-break,normal); overflow-wrap: anywhere; }

.VfPpkd-suEOdc-OWXEXe-eo9XGd-RCfa3e .VfPpkd-z59Tgd-OiiCO { transition: opacity 0.15s cubic-bezier(0, 0, 0.2, 1) 0ms, transform 0.15s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.15s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-suEOdc-OWXEXe-ZYIfFd-RCfa3e .VfPpkd-z59Tgd-OiiCO { transition: opacity 75ms cubic-bezier(0.4, 0, 1, 1) 0ms; }

.VfPpkd-suEOdc { position: fixed; display: none; z-index: 9; }

.VfPpkd-suEOdc-sM5MNb-OWXEXe-nzrxxc { position: relative; }

.VfPpkd-suEOdc-OWXEXe-TSZdd, .VfPpkd-suEOdc-OWXEXe-eo9XGd, .VfPpkd-suEOdc-OWXEXe-ZYIfFd { display: inline-flex; }

.VfPpkd-suEOdc-OWXEXe-TSZdd.VfPpkd-suEOdc-OWXEXe-nzrxxc, .VfPpkd-suEOdc-OWXEXe-eo9XGd.VfPpkd-suEOdc-OWXEXe-nzrxxc, .VfPpkd-suEOdc-OWXEXe-ZYIfFd.VfPpkd-suEOdc-OWXEXe-nzrxxc { display: inline-block; left: -320px; position: absolute; }

.VfPpkd-z59Tgd { line-height: 16px; padding: 4px 8px; min-width: 40px; max-width: 200px; min-height: 24px; max-height: 40vh; box-sizing: border-box; overflow: hidden; text-align: center; }

.VfPpkd-z59Tgd::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 1px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-z59Tgd::before { border-color: canvastext; }
}

.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd { -webkit-box-align: start; align-items: flex-start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; min-height: 24px; min-width: 40px; max-width: 320px; position: relative; }

.VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd { text-align: left; }

[dir="rtl"] .VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd, .VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd[dir="rtl"] { text-align: right; }

.VfPpkd-z59Tgd .VfPpkd-MlC99b { margin: 0px 8px; }

.VfPpkd-z59Tgd .VfPpkd-IqDDtd { max-width: 184px; margin: 8px; text-align: left; }

[dir="rtl"] .VfPpkd-z59Tgd .VfPpkd-IqDDtd, .VfPpkd-z59Tgd .VfPpkd-IqDDtd[dir="rtl"] { text-align: right; }

.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-IqDDtd { max-width: 304px; align-self: stretch; }

.VfPpkd-z59Tgd .VfPpkd-IqDDtd-hSRGPd { text-decoration: none; }

.VfPpkd-suEOdc-OWXEXe-nzrxxc-LQLjdd, .VfPpkd-IqDDtd, .VfPpkd-MlC99b { z-index: 1; }

.VfPpkd-z59Tgd-OiiCO { opacity: 0; transform: scale(0.8); will-change: transform, opacity; }

.VfPpkd-suEOdc-OWXEXe-TSZdd .VfPpkd-z59Tgd-OiiCO { transform: scale(1); opacity: 1; }

.VfPpkd-suEOdc-OWXEXe-ZYIfFd .VfPpkd-z59Tgd-OiiCO { transform: scale(1); }

.VfPpkd-Djsh7e-XxIAqe-ma6Yeb, .VfPpkd-Djsh7e-XxIAqe-cGMI2b { position: absolute; height: 24px; width: 24px; transform: rotate(35deg) skewY(20deg) scaleX(0.939693); }

.VfPpkd-Djsh7e-XxIAqe-ma6Yeb .VfPpkd-BFbNVe-bF1uUb, .VfPpkd-Djsh7e-XxIAqe-cGMI2b .VfPpkd-BFbNVe-bF1uUb { width: 100%; height: 100%; top: 0px; left: 0px; }

.VfPpkd-Djsh7e-XxIAqe-cGMI2b { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 1px -2px, rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 1px 5px 0px; outline: transparent solid 1px; z-index: -1; }

@media screen and (forced-colors: active) {
  .VfPpkd-Djsh7e-XxIAqe-cGMI2b { outline-color: canvastext; }
}

.VfPpkd-BFbNVe-bF1uUb { position: absolute; border-radius: inherit; pointer-events: none; opacity: var(--mdc-elevation-overlay-opacity,0); transition: opacity 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; background-color: var(--mdc-elevation-overlay-color,#fff); }

.NZp2ef { background-color: rgb(232, 234, 237); }

.EY8ABd { z-index: 2101; }

.EY8ABd .VfPpkd-z59Tgd { background-color: rgb(60, 64, 67); color: rgb(232, 234, 237); }

.EY8ABd .VfPpkd-MlC99b, .EY8ABd .VfPpkd-IqDDtd { color: rgb(60, 64, 67); }

.EY8ABd .VfPpkd-IqDDtd-hSRGPd { color: rgb(26, 115, 232); }

.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd, .EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb, .EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b { background-color: rgb(255, 255, 255); }

.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; }

.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd { border-radius: 8px; }

.ziykHb { z-index: 2101; }

.ziykHb .VfPpkd-z59Tgd { background-color: rgb(60, 64, 67); color: rgb(232, 234, 237); }

.ziykHb .VfPpkd-MlC99b, .ziykHb .VfPpkd-IqDDtd { color: rgb(60, 64, 67); }

.ziykHb .VfPpkd-IqDDtd-hSRGPd { color: rgb(26, 115, 232); }

.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd, .ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb, .ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b { background-color: rgb(255, 255, 255); }

.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; }

.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd { border-radius: 8px; }

.EY8ABd-OWXEXe-TAWMXe { position: absolute; left: -10000px; top: auto; width: 1px; height: 1px; overflow: hidden; user-select: none; }

@-webkit-keyframes mdc-ripple-fg-radius-in { 
  0% { animation-timing-function: cubic-bezier(0.4, 0, 0.2, 1); transform: translate(var(--mdc-ripple-fg-translate-start,0)) scale(1); }
  100% { transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }
}

@keyframes mdc-ripple-fg-radius-in { 
  0% { animation-timing-function: cubic-bezier(0.4, 0, 0.2, 1); transform: translate(var(--mdc-ripple-fg-translate-start,0)) scale(1); }
  100% { transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }
}

@-webkit-keyframes mdc-ripple-fg-opacity-in { 
  0% { animation-timing-function: linear; opacity: 0; }
  100% { opacity: var(--mdc-ripple-fg-opacity,0); }
}

@keyframes mdc-ripple-fg-opacity-in { 
  0% { animation-timing-function: linear; opacity: 0; }
  100% { opacity: var(--mdc-ripple-fg-opacity,0); }
}

@-webkit-keyframes mdc-ripple-fg-opacity-out { 
  0% { animation-timing-function: linear; opacity: var(--mdc-ripple-fg-opacity,0); }
  100% { opacity: 0; }
}

@keyframes mdc-ripple-fg-opacity-out { 
  0% { animation-timing-function: linear; opacity: var(--mdc-ripple-fg-opacity,0); }
  100% { opacity: 0; }
}

.VfPpkd-ksKsZd-XxIAqe { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; position: relative; outline: none; overflow: hidden; }

.VfPpkd-ksKsZd-XxIAqe::before, .VfPpkd-ksKsZd-XxIAqe::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-ksKsZd-XxIAqe::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-ksKsZd-XxIAqe::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf::after { animation: 150ms ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-ksKsZd-XxIAqe::before, .VfPpkd-ksKsZd-XxIAqe::after { top: calc(-50%); left: calc(-50%); width: 200%; height: 200%; }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded], .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd { overflow: visible; }

.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::before, .VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::after, .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::before, .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after { top: calc(0%); left: calc(0%); width: 100%; height: 100%; }

.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::before, .VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after, .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::before, .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after { top: var(--mdc-ripple-top,calc(50% - 50%)); left: var(--mdc-ripple-left,calc(50% - 50%)); width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after, .VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-ksKsZd-XxIAqe::before, .VfPpkd-ksKsZd-XxIAqe::after { background-color: var(--mdc-ripple-color,#000); }

.VfPpkd-ksKsZd-XxIAqe:hover::before, .VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE::before { opacity: var(--mdc-ripple-hover-opacity,0.04); }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before, .VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):focus::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0.12); }

.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d)::after { transition: opacity 150ms linear 0s; }

.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):active::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-Bz112c-LgbsSe { font-size: 24px; width: 48px; height: 48px; padding: 12px; }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 48px; max-width: 48px; }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 40px; height: 40px; margin: 4px; }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 40px; max-width: 40px; }

.VfPpkd-Bz112c-LgbsSe:disabled { color: var(--mdc-theme-text-disabled-on-light,rgba(0,0,0,.38)); }

.VfPpkd-Bz112c-LgbsSe svg, .VfPpkd-Bz112c-LgbsSe img { width: 24px; height: 24px; }

.VfPpkd-Bz112c-LgbsSe { display: inline-block; position: relative; box-sizing: border-box; border: none; outline: none; background-color: transparent; fill: currentcolor; color: inherit; text-decoration: none; cursor: pointer; user-select: none; z-index: 0; overflow: visible; }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 48px; left: 50%; width: 48px; transform: translate(-50%, -50%); }

@media screen and (forced-colors: active) {
  .VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-J1Ukfc-LhBDec, .VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-J1Ukfc-LhBDec { display: block; }
}

.VfPpkd-Bz112c-LgbsSe:disabled { cursor: default; pointer-events: none; }

.VfPpkd-Bz112c-LgbsSe[hidden] { display: none; }

.VfPpkd-Bz112c-LgbsSe-OWXEXe-KVuj8d-Q3DXx { -webkit-box-align: center; align-items: center; display: inline-flex; -webkit-box-pack: center; justify-content: center; }

.VfPpkd-Bz112c-J1Ukfc-LhBDec { pointer-events: none; border: 2px solid transparent; border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: 100%; width: 100%; display: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-Bz112c-J1Ukfc-LhBDec { border-color: canvastext; }
}

.VfPpkd-Bz112c-J1Ukfc-LhBDec::after { content: ""; border: 2px solid transparent; border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .VfPpkd-Bz112c-J1Ukfc-LhBDec::after { border-color: canvastext; }
}

.VfPpkd-Bz112c-kBDsod { display: inline-block; }

.VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd, .VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod { display: none; }

.VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd { display: inline-block; }

.VfPpkd-Bz112c-mRLv6 { height: 100%; left: 0px; outline: none; position: absolute; top: 0px; width: 100%; }

.VfPpkd-Bz112c-LgbsSe { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Bz112c-Jh9lGc::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Bz112c-Jh9lGc::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Bz112c-Jh9lGc::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after { top: 0px; left: 0px; width: 100%; height: 100%; }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after { background-color: var(--mdc-ripple-color,#000); }

.VfPpkd-Bz112c-LgbsSe:hover .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-Bz112c-LgbsSe:disabled:hover .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before, .VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc { height: 100%; left: 0px; pointer-events: none; position: absolute; top: 0px; width: 100%; z-index: -1; }

.VfPpkd-dgl2Hf-ppHlrf-sM5MNb { display: inline; }

.VfPpkd-LgbsSe { position: relative; display: inline-flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; box-sizing: border-box; min-width: 64px; border: none; outline: none; line-height: inherit; user-select: none; appearance: none; overflow: visible; vertical-align: middle; background: transparent; }

.VfPpkd-LgbsSe .VfPpkd-BFbNVe-bF1uUb { width: 100%; height: 100%; top: 0px; left: 0px; }

.VfPpkd-LgbsSe:active { outline: none; }

.VfPpkd-LgbsSe:hover { cursor: pointer; }

.VfPpkd-LgbsSe:disabled { cursor: default; pointer-events: none; }

.VfPpkd-LgbsSe[hidden] { display: none; }

.VfPpkd-LgbsSe .VfPpkd-kBDsod { margin-left: 0px; margin-right: 8px; display: inline-block; position: relative; vertical-align: top; }

[dir="rtl"] .VfPpkd-LgbsSe .VfPpkd-kBDsod, .VfPpkd-LgbsSe .VfPpkd-kBDsod[dir="rtl"] { margin-left: 8px; margin-right: 0px; }

.VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge { font-size: 0px; position: absolute; transform: translate(-50%, -50%); top: 50%; left: 50%; line-height: normal; }

.VfPpkd-LgbsSe .VfPpkd-vQzf8d { position: relative; }

.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec { pointer-events: none; border: 2px solid transparent; border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); display: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec { border-color: canvastext; }
}

.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after { content: ""; border: 2px solid transparent; border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after { border-color: canvastext; }
}

@media screen and (forced-colors: active) {
  .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-J1Ukfc-LhBDec, .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-J1Ukfc-LhBDec { display: block; }
}

.VfPpkd-LgbsSe .VfPpkd-RLmnJb { position: absolute; top: 50%; height: 48px; left: 0px; right: 0px; transform: translateY(-50%); }

.VfPpkd-vQzf8d + .VfPpkd-kBDsod { margin-left: 8px; margin-right: 0px; }

[dir="rtl"] .VfPpkd-vQzf8d + .VfPpkd-kBDsod, .VfPpkd-vQzf8d + .VfPpkd-kBDsod[dir="rtl"] { margin-left: 0px; margin-right: 8px; }

svg.VfPpkd-kBDsod { fill: currentcolor; }

.VfPpkd-LgbsSe-OWXEXe-dgl2Hf { margin-top: 6px; margin-bottom: 6px; }

.VfPpkd-LgbsSe { -webkit-font-smoothing: antialiased; text-decoration: none; }

.VfPpkd-LgbsSe { padding: 0px 8px; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ { transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; padding: 0px 16px; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 12px 0px 16px; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 16px 0px 12px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb { transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; padding: 0px 16px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 12px 0px 16px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 16px 0px 12px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc { border-style: solid; transition: border 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc { border-style: solid; border-color: transparent; }

.VfPpkd-LgbsSe { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: 1; }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after { z-index: 0; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Jh9lGc::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Jh9lGc::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Jh9lGc::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after { top: -50%; left: -50%; width: 200%; height: 200%; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-Jh9lGc { position: absolute; box-sizing: content-box; overflow: hidden; z-index: 0; inset: 0px; }

.VfPpkd-LgbsSe { font-family: Roboto, sans-serif; font-size: 0.875rem; letter-spacing: 0.0892857em; font-weight: 500; text-transform: uppercase; height: 36px; border-radius: 4px; }

.VfPpkd-LgbsSe:not(:disabled) { color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe:disabled { color: rgba(0, 0, 0, 0.38); }

.VfPpkd-LgbsSe .VfPpkd-kBDsod { font-size: 1.125rem; width: 1.125rem; height: 1.125rem; }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after { background-color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: 0.04; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: 0.12; }

.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: 0.12; }

.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-text-button-pressed-state-layer-opacity,0.12); }

.VfPpkd-LgbsSe .VfPpkd-Jh9lGc { border-radius: 4px; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ { font-family: Roboto, sans-serif; font-size: 0.875rem; letter-spacing: 0.0892857em; font-weight: 500; text-transform: uppercase; height: 36px; border-radius: 4px; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled) { background-color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled { background-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled) { color: rgb(255, 255, 255); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled { color: rgba(0, 0, 0, 0.38); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-kBDsod { font-size: 1.125rem; width: 1.125rem; height: 1.125rem; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::after { background-color: rgb(255, 255, 255); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:hover .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: 0.08; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: 0.24; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: 0.24; }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-filled-button-pressed-state-layer-opacity,0.24); }

.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc { border-radius: 4px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb { font-family: Roboto, sans-serif; font-size: 0.875rem; letter-spacing: 0.0892857em; font-weight: 500; text-transform: uppercase; height: 36px; border-radius: 4px; box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 1px -2px, rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 1px 5px 0px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled) { background-color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled { background-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled) { color: rgb(255, 255, 255); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled { color: rgba(0, 0, 0, 0.38); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-kBDsod { font-size: 1.125rem; width: 1.125rem; height: 1.125rem; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::after { background-color: rgb(255, 255, 255); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: 0.08; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: 0.24; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: 0.24; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-protected-button-pressed-state-layer-opacity,0.24); }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc { border-radius: 4px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus { box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px -1px, rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover { box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px -1px, rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled):active { box-shadow: rgba(0, 0, 0, 0.2) 0px 5px 5px -3px, rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px; }

.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled { box-shadow: rgba(0, 0, 0, 0.2) 0px 0px 0px 0px, rgba(0, 0, 0, 0.14) 0px 0px 0px 0px, rgba(0, 0, 0, 0.12) 0px 0px 0px 0px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc { font-family: Roboto, sans-serif; font-size: 0.875rem; letter-spacing: 0.0892857em; font-weight: 500; text-transform: uppercase; height: 36px; border-radius: 4px; padding: 0px 15px; border-width: 1px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled) { color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled { color: rgba(0, 0, 0, 0.38); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-kBDsod { font-size: 1.125rem; width: 1.125rem; height: 1.125rem; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::after { background-color: rgb(98, 0, 238); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:hover .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: 0.04; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: 0.12; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: 0.12; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-outlined-button-pressed-state-layer-opacity,0.12); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc { border-radius: 4px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled) { border-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled { border-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 11px 0px 15px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 15px 0px 11px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc { inset: -1px; border-width: 1px; }

.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-RLmnJb { left: -1px; width: calc(100% + 2px); }

.nCP5yc { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; transition: border 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s, box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; box-shadow: none; }

.nCP5yc .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.nCP5yc:not(:disabled) { background-color: var(--gm-fillbutton-container-color,rgb(26,115,232)); }

.nCP5yc:not(:disabled) { color: var(--gm-fillbutton-ink-color,#fff); }

.nCP5yc:disabled { background-color: var(--gm-fillbutton-disabled-container-color,rgba(60,64,67,.12)); }

.nCP5yc:disabled { color: var(--gm-fillbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.nCP5yc .VfPpkd-Jh9lGc::before, .nCP5yc .VfPpkd-Jh9lGc::after { background-color: var(--gm-fillbutton-state-color,rgb(32,33,36)); }

.nCP5yc:hover .VfPpkd-Jh9lGc::before, .nCP5yc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.16); }

.nCP5yc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.24); }

.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.2); }

.nCP5yc.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.2); }

.nCP5yc .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(255, 255, 255); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.nCP5yc:hover { box-shadow: 0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.nCP5yc:hover .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.nCP5yc:active { box-shadow: 0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.nCP5yc:active .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.nCP5yc:disabled { box-shadow: none; }

.nCP5yc:disabled:hover .VfPpkd-Jh9lGc::before, .nCP5yc:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.nCP5yc:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.nCP5yc:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.nCP5yc:disabled .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Rj2Mlf { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; transition: border 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s, box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; box-shadow: none; }

.Rj2Mlf .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.Rj2Mlf:not(:disabled) { color: var(--gm-hairlinebutton-ink-color,rgb(26,115,232)); }

.Rj2Mlf:not(:disabled) { border-color: var(--gm-hairlinebutton-outline-color,rgb(218,220,224)); }

.Rj2Mlf:not(:disabled):hover { border-color: var(--gm-hairlinebutton-outline-color,rgb(218,220,224)); }

.Rj2Mlf:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .Rj2Mlf:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus { border-color: var(--gm-hairlinebutton-outline-color--stateful,rgb(23,78,166)); }

.Rj2Mlf:not(:disabled):active, .Rj2Mlf:not(:disabled):focus:active { border-color: var(--gm-hairlinebutton-outline-color,rgb(218,220,224)); }

.Rj2Mlf:disabled { color: var(--gm-hairlinebutton-disabled-ink-color,rgba(60,64,67,.38)); }

.Rj2Mlf:disabled { border-color: var(--gm-hairlinebutton-disabled-outline-color,rgba(60,64,67,.12)); }

.Rj2Mlf:hover:not(:disabled), .Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled), .Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled), .Rj2Mlf:active:not(:disabled) { color: var(--gm-hairlinebutton-ink-color--stateful,rgb(23,78,166)); }

.Rj2Mlf .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(26, 115, 232); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.Rj2Mlf .VfPpkd-Jh9lGc::before, .Rj2Mlf .VfPpkd-Jh9lGc::after { background-color: var(--gm-hairlinebutton-state-color,rgb(26,115,232)); }

.Rj2Mlf:hover .VfPpkd-Jh9lGc::before, .Rj2Mlf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.Rj2Mlf:disabled:hover .VfPpkd-Jh9lGc::before, .Rj2Mlf:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.Rj2Mlf:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.Rj2Mlf:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.b9hyVd { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; transition: border 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s, box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; border-width: 0px; box-shadow: 0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.b9hyVd .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.b9hyVd:not(:disabled) { background-color: var(--gm-protectedbutton-container-color,#fff); }

.b9hyVd:not(:disabled) { color: var(--gm-protectedbutton-ink-color,rgb(26,115,232)); }

.b9hyVd:disabled { background-color: var(--gm-protectedbutton-disabled-container-color,rgba(60,64,67,.12)); }

.b9hyVd:disabled { color: var(--gm-protectedbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.b9hyVd:hover:not(:disabled), .b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled), .b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled), .b9hyVd:active:not(:disabled) { color: var(--gm-protectedbutton-ink-color--stateful,rgb(23,78,166)); }

.b9hyVd .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(26, 115, 232); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus { border-width: 0px; box-shadow: 0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-BFbNVe-bF1uUb, .b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.b9hyVd:hover { border-width: 0px; box-shadow: 0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.b9hyVd:hover .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.b9hyVd:not(:disabled):active { border-width: 0px; box-shadow: 0 1px 3px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 4px 8px 3px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15)); }

.b9hyVd:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.b9hyVd .VfPpkd-Jh9lGc::before, .b9hyVd .VfPpkd-Jh9lGc::after { background-color: var(--gm-protectedbutton-state-color,rgb(26,115,232)); }

.b9hyVd:hover .VfPpkd-Jh9lGc::before, .b9hyVd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.b9hyVd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.b9hyVd:disabled { box-shadow: none; }

.b9hyVd:disabled .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.b9hyVd:disabled:hover .VfPpkd-Jh9lGc::before, .b9hyVd:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.b9hyVd:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.b9hyVd:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.Kjnxrf { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; transition: border 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s, box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; box-shadow: none; }

.Kjnxrf .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.Kjnxrf:not(:disabled) { background-color: rgb(232, 240, 254); }

.Kjnxrf:not(:disabled) { color: rgb(25, 103, 210); }

.Kjnxrf:disabled { background-color: rgba(60, 64, 67, 0.12); }

.Kjnxrf:disabled { color: rgba(60, 64, 67, 0.38); }

.Kjnxrf:hover:not(:disabled), .Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled), .Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled), .Kjnxrf:active:not(:disabled) { color: rgb(23, 78, 166); }

.Kjnxrf .VfPpkd-Jh9lGc::before, .Kjnxrf .VfPpkd-Jh9lGc::after { background-color: var(--mdc-ripple-color,rgb(25,103,210)); }

.Kjnxrf:hover .VfPpkd-Jh9lGc::before, .Kjnxrf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.Kjnxrf.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.Kjnxrf .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(25, 103, 210); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.Kjnxrf:hover { box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.Kjnxrf:hover .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Kjnxrf:not(:disabled):active { box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.Kjnxrf:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Kjnxrf:disabled { box-shadow: none; }

.Kjnxrf:disabled .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.Kjnxrf:disabled:hover .VfPpkd-Jh9lGc::before, .Kjnxrf:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.Kjnxrf:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.Kjnxrf:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.ksBjEc { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; }

.ksBjEc .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.ksBjEc:not(:disabled) { background-color: transparent; }

.ksBjEc:not(:disabled) { color: var(--gm-colortextbutton-ink-color,rgb(26,115,232)); }

.ksBjEc:disabled { color: var(--gm-colortextbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(26, 115, 232); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.ksBjEc:hover:not(:disabled), .ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled), .ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled), .ksBjEc:active:not(:disabled) { color: var(--gm-colortextbutton-ink-color--stateful,rgb(23,78,166)); }

.ksBjEc .VfPpkd-Jh9lGc::before, .ksBjEc .VfPpkd-Jh9lGc::after { background-color: var(--gm-colortextbutton-state-color,rgb(26,115,232)); }

.ksBjEc:hover .VfPpkd-Jh9lGc::before, .ksBjEc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.ksBjEc.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.ksBjEc:disabled:hover .VfPpkd-Jh9lGc::before, .ksBjEc:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.ksBjEc:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.ksBjEc:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.LjDxcd { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0107143em; font-weight: 500; text-transform: none; }

.LjDxcd .VfPpkd-Jh9lGc { height: 100%; position: absolute; overflow: hidden; width: 100%; z-index: 0; }

.LjDxcd:not(:disabled) { color: var(--gm-neutraltextbutton-ink-color,rgb(95,99,104)); }

.LjDxcd:disabled { color: var(--gm-neutraltextbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.LjDxcd:hover:not(:disabled), .LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled), .LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled), .LjDxcd:active:not(:disabled) { color: var(--gm-neutraltextbutton-ink-color--stateful,rgb(32,33,36)); }

.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(95, 99, 104); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo, .LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.LjDxcd .VfPpkd-Jh9lGc::before, .LjDxcd .VfPpkd-Jh9lGc::after { background-color: var(--gm-neutraltextbutton-state-color,rgb(95,99,104)); }

.LjDxcd:hover .VfPpkd-Jh9lGc::before, .LjDxcd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.LjDxcd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.LjDxcd:disabled:hover .VfPpkd-Jh9lGc::before, .LjDxcd:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before { opacity: var(--mdc-ripple-hover-opacity,0); }

.LjDxcd:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before, .LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,0); }

.LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after { transition: opacity 0.15s linear 0s; }

.LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,0); }

.LjDxcd:disabled.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0); }

.DuMIQc { padding: 0px 24px; }

.P62QJc { padding: 0px 23px; border-width: 1px; }

.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 11px 0px 23px; }

.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 23px 0px 11px; }

.P62QJc .VfPpkd-Jh9lGc { inset: -1px; border-width: 1px; }

.P62QJc .VfPpkd-RLmnJb { left: -1px; width: calc(100% + 2px); }

.yHy1rc { z-index: 0; }

.yHy1rc .VfPpkd-Bz112c-Jh9lGc::before, .yHy1rc .VfPpkd-Bz112c-Jh9lGc::after { z-index: -1; }

.yHy1rc:disabled { color: var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.fzRBVc { z-index: 0; }

.fzRBVc .VfPpkd-Bz112c-Jh9lGc::before, .fzRBVc .VfPpkd-Bz112c-Jh9lGc::after { z-index: -1; }

.fzRBVc:disabled { color: var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38)); }

.WpHeLc { height: 100%; left: 0px; position: absolute; top: 0px; width: 100%; outline: none; }

[dir="rtl"] .HDnnrf .VfPpkd-kBDsod, .HDnnrf .VfPpkd-kBDsod[dir="rtl"] { transform: scaleX(-1); }

[dir="rtl"] .QDwDD, .QDwDD[dir="rtl"] { transform: scaleX(-1); }

.PDpWxe { will-change: unset; }

.LQeN7 .VfPpkd-J1Ukfc-LhBDec { pointer-events: none; border: 2px solid rgb(24, 90, 188); border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .LQeN7 .VfPpkd-J1Ukfc-LhBDec { border-color: canvastext; }
}

.LQeN7 .VfPpkd-J1Ukfc-LhBDec::after { content: ""; border: 2px solid rgb(232, 240, 254); border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .LQeN7 .VfPpkd-J1Ukfc-LhBDec::after { border-color: canvastext; }
}

.LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec { display: inline-block; }

@media (-ms-high-contrast:active), (-ms-high-contrast:none) {
  .LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec { display: none; }
}

.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec { pointer-events: none; border: 2px solid rgb(24, 90, 188); border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: 100%; width: 100%; }

@media screen and (forced-colors: active) {
  .mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec { border-color: canvastext; }
}

.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after { content: ""; border: 2px solid rgb(232, 240, 254); border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after { border-color: canvastext; }
}

.mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec { display: inline-block; }

@media (-ms-high-contrast:active), (-ms-high-contrast:none) {
  .mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec { display: none; }
}

.MyRpB .VfPpkd-kBDsod, .MyRpB .VfPpkd-vQzf8d { opacity: 0; }

[data-tooltip-enabled="true"]:disabled, .VfPpkd-Bz112c-LgbsSe[data-tooltip-enabled="true"]:disabled .VfPpkd-Bz112c-Jh9lGc { pointer-events: auto; }

.xFWpbf { border-radius: var(--dt-corner-button,.25rem); }

.xFWpbf::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 1px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .xFWpbf::before { border-color: canvastext; }
}

.vhoiae .xFWpbf, .X9XeLb .xFWpbf, .cWKK1c .xFWpbf, .aJfoSc .xFWpbf, .TOb6Ze .xFWpbf { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,.0178571429em); text-overflow: ellipsis; white-space: nowrap; }

.xFWpbf .VfPpkd-Jh9lGc { border-radius: inherit; }

.xFWpbf:disabled { color: var(--dt-on-disabled,rgba(60,64,67,.38)); }

.uJtSke.kphldf { --gm-hairlinebutton-outline-color: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-outline-color--stateful: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-ink-color: var(--dt-error-action,rgb(197,34,31)); --gm-hairlinebutton-ink-color--stateful: var(--dt-error-action-stateful,rgb(179,20,18)); --gm-hairlinebutton-state-color: var(--dt-error-action-state-layer,rgb(197,34,31)); }

.uJtSke.rNe0id { --gm-hairlinebutton-outline-color: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-outline-color--stateful: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-ink-color: var(--dt-warning-action,rgb(60,64,67)); --gm-hairlinebutton-ink-color--stateful: var(--dt-warning-action-stateful,rgb(32,33,36)); --gm-hairlinebutton-state-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); }

.uJtSke.sj692e { --gm-hairlinebutton-outline-color: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-outline-color--stateful: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-hairlinebutton-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); --gm-hairlinebutton-state-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); }

.uJtSke.IY5c4e { --gm-hairlinebutton-outline-color: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-outline-color--stateful: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-ink-color: var(--dt-tertiary-action,rgb(19,115,51)); --gm-hairlinebutton-ink-color--stateful: var(--dt-tertiary-action-stateful,rgb(13,101,45)); --gm-hairlinebutton-state-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); }

.uJtSke.qoCZef { --gm-hairlinebutton-outline-color: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-outline-color--stateful: var(--dt-outline,rgb(128,134,139)); --gm-hairlinebutton-ink-color: var(--dt-neutral-action,rgb(60,64,67)); --gm-hairlinebutton-ink-color--stateful: var(--dt-neutral-action-stateful,rgb(32,33,36)); --gm-hairlinebutton-state-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); }

.uJtSke:disabled { border-color: var(--dt-disabled,rgba(60,64,67,.12)); }

.oWBWHf.kphldf { --gm-fillbutton-container-color: var(--dt-error,rgb(217,48,37)); --gm-fillbutton-ink-color: var(--dt-on-error,#fff); --gm-fillbutton-state-color: var(--dt-inverse-surface,rgb(32,33,36)); }

.oWBWHf.rNe0id { --gm-fillbutton-container-color: var(--dt-warning,rgb(249,171,0)); --gm-fillbutton-ink-color: var(--dt-on-warning,rgb(32,33,36)); --gm-fillbutton-state-color: var(--dt-inverse-surface,rgb(32,33,36)); }

.oWBWHf.sj692e { --gm-fillbutton-container-color: var(--dt-primary,rgb(26,115,232)); --gm-fillbutton-ink-color: var(--dt-on-primary,#fff); --gm-fillbutton-state-color: var(--dt-inverse-surface,rgb(32,33,36)); }

.oWBWHf.IY5c4e { --gm-fillbutton-container-color: var(--dt-tertiary,rgb(24,128,56)); --gm-fillbutton-ink-color: var(--dt-on-tertiary,#fff); --gm-fillbutton-state-color: var(--dt-inverse-surface,rgb(32,33,36)); }

.oWBWHf.qoCZef { --gm-fillbutton-container-color: var(--dt-neutral,rgb(60,64,67)); --gm-fillbutton-ink-color: var(--dt-on-neutral,#fff); --gm-fillbutton-state-color: var(--dt-inverse-surface,rgb(32,33,36)); }

.oWBWHf:disabled { background-color: var(--dt-disabled,rgba(60,64,67,.12)); }

.hLvULc.kphldf { --gm-protectedbutton-container-color: var(--dt-background,#fff); --gm-protectedbutton-ink-color: var(--dt-error-action,rgb(197,34,31)); --gm-protectedbutton-ink-color--stateful: var(--dt-error-action-stateful,rgb(179,20,18)); --gm-protectedbutton-state-color: var(--dt-error-action-state-layer,rgb(197,34,31)); }

.hLvULc.rNe0id { --gm-protectedbutton-container-color: var(--dt-background,#fff); --gm-protectedbutton-ink-color: var(--dt-warning-action,rgb(60,64,67)); --gm-protectedbutton-ink-color--stateful: var(--dt-warning-action-stateful,rgb(32,33,36)); --gm-protectedbutton-state-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); }

.hLvULc.sj692e { --gm-protectedbutton-container-color: var(--dt-background,#fff); --gm-protectedbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-protectedbutton-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); --gm-protectedbutton-state-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); }

.hLvULc.IY5c4e { --gm-protectedbutton-container-color: var(--dt-background,#fff); --gm-protectedbutton-ink-color: var(--dt-tertiary-action,rgb(19,115,51)); --gm-protectedbutton-ink-color--stateful: var(--dt-tertiary-action-stateful,rgb(13,101,45)); --gm-protectedbutton-state-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); }

.hLvULc.qoCZef { --gm-protectedbutton-container-color: var(--dt-background,#fff); --gm-protectedbutton-ink-color: var(--dt-neutral-action,rgb(60,64,67)); --gm-protectedbutton-ink-color--stateful: var(--dt-neutral-action-stateful,rgb(32,33,36)); --gm-protectedbutton-state-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); }

.vhoiae .uFAPIe, .X9XeLb .uFAPIe, .cWKK1c .uFAPIe, .aJfoSc .uFAPIe, .TOb6Ze .uFAPIe { padding: 0px 12px; border-width: 1px; }

.vhoiae .uFAPIe:not(:disabled), .X9XeLb .uFAPIe:not(:disabled), .cWKK1c .uFAPIe:not(:disabled), .aJfoSc .uFAPIe:not(:disabled), .TOb6Ze .uFAPIe:not(:disabled) { border-color: transparent; }

.vhoiae .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .X9XeLb .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .cWKK1c .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .aJfoSc .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .TOb6Ze .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 11px 0px 12px; }

.vhoiae .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .X9XeLb .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .cWKK1c .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .aJfoSc .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .TOb6Ze .uFAPIe.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 12px 0px 11px; }

.vhoiae .uFAPIe .VfPpkd-Jh9lGc, .X9XeLb .uFAPIe .VfPpkd-Jh9lGc, .cWKK1c .uFAPIe .VfPpkd-Jh9lGc, .aJfoSc .uFAPIe .VfPpkd-Jh9lGc, .TOb6Ze .uFAPIe .VfPpkd-Jh9lGc { inset: -1px; border-width: 1px; }

.vhoiae .uFAPIe .VfPpkd-RLmnJb, .X9XeLb .uFAPIe .VfPpkd-RLmnJb, .cWKK1c .uFAPIe .VfPpkd-RLmnJb, .aJfoSc .uFAPIe .VfPpkd-RLmnJb, .TOb6Ze .uFAPIe .VfPpkd-RLmnJb { left: -1px; width: calc(100% + 2px); }

.vhoiae .uFAPIe.cd29Sd, .X9XeLb .uFAPIe.cd29Sd, .cWKK1c .uFAPIe.cd29Sd, .aJfoSc .uFAPIe.cd29Sd, .TOb6Ze .uFAPIe.cd29Sd { padding-right: 16px; }

.uFAPIe.kphldf { --gm-colortextbutton-ink-color: var(--dt-error-action,rgb(197,34,31)); --gm-colortextbutton-state-color: var(--dt-error-action-state-layer,rgb(197,34,31)); --gm-colortextbutton-ink-color--stateful: var(--dt-error-action-stateful,rgb(179,20,18)); }

.uFAPIe.rNe0id { --gm-colortextbutton-ink-color: var(--dt-warning-action,rgb(60,64,67)); --gm-colortextbutton-state-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); --gm-colortextbutton-ink-color--stateful: var(--dt-warning-action-stateful,rgb(32,33,36)); }

.uFAPIe.sj692e { --gm-colortextbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-colortextbutton-state-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); --gm-colortextbutton-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); }

.uFAPIe.IY5c4e { --gm-colortextbutton-ink-color: var(--dt-tertiary-action,rgb(19,115,51)); --gm-colortextbutton-state-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); --gm-colortextbutton-ink-color--stateful: var(--dt-tertiary-action-stateful,rgb(13,101,45)); }

.uFAPIe.qoCZef { --gm-colortextbutton-ink-color: var(--dt-neutral-action,rgb(60,64,67)); --gm-colortextbutton-state-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); --gm-colortextbutton-ink-color--stateful: var(--dt-neutral-action-stateful,rgb(32,33,36)); }

.uFAPIe.bustDd.sj692e { --gm-colortextbutton-ink-color: var(--dt-on-primary,#fff); --gm-colortextbutton-state-color: var(--dt-on-primary,#fff); --gm-colortextbutton-ink-color--stateful: var(--dt-on-primary,#fff); }

.uFAPIe.bustDd.IY5c4e { --gm-colortextbutton-ink-color: var(--dt-on-tertiary,#fff); --gm-colortextbutton-state-color: var(--dt-on-tertiary,#fff); --gm-colortextbutton-ink-color--stateful: var(--dt-on-tertiary,#fff); }

.uFAPIe.bustDd.qoCZef { --gm-colortextbutton-ink-color: var(--dt-on-neutral,#fff); --gm-colortextbutton-state-color: var(--dt-on-neutral,#fff); --gm-colortextbutton-ink-color--stateful: var(--dt-on-neutral,#fff); }

.uFAPIe.bustDd.kphldf { --gm-colortextbutton-ink-color: var(--dt-on-error,#fff); --gm-colortextbutton-state-color: var(--dt-on-error,#fff); --gm-colortextbutton-ink-color--stateful: var(--dt-on-error,#fff); }

.uFAPIe.bustDd.rNe0id { --gm-colortextbutton-ink-color: var(--dt-on-warning,rgb(32,33,36)); --gm-colortextbutton-state-color: var(--dt-on-warning,rgb(32,33,36)); --gm-colortextbutton-ink-color--stateful: var(--dt-on-warning,rgb(32,33,36)); }

.p9NqC { border-width: 1px; padding: 12px; }

.p9NqC:not(:disabled) { border-color: transparent; }

.p9NqC.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 11px 0px 12px; }

.p9NqC.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 12px 0px 11px; }

.p9NqC .VfPpkd-Jh9lGc { inset: -1px; border-width: 1px; }

.p9NqC .VfPpkd-RLmnJb { left: -1px; width: calc(100% + 2px); }

.p9NqC:focus, .p9NqC:hover, .p9NqC:active { border-width: 2px; padding: 12px; outline: transparent solid 2px; }

.p9NqC:focus.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .p9NqC:hover.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg, .p9NqC:active.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg { padding: 0px 10px 0px 12px; }

.p9NqC:focus.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .p9NqC:hover.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc, .p9NqC:active.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc { padding: 0px 12px 0px 10px; }

.p9NqC:focus .VfPpkd-Jh9lGc, .p9NqC:hover .VfPpkd-Jh9lGc, .p9NqC:active .VfPpkd-Jh9lGc { inset: -2px; border-width: 2px; }

.p9NqC:focus .VfPpkd-RLmnJb, .p9NqC:hover .VfPpkd-RLmnJb, .p9NqC:active .VfPpkd-RLmnJb { left: -2px; width: calc(100% + 4px); }

.p9NqC.kphldf { --mdc-ripple-color: var(--dt-error-action-state-layer,rgb(197,34,31)); --gm-iconbutton-ink-color: var(--dt-error-action,rgb(197,34,31)); }

.p9NqC.kphldf:focus, .p9NqC.kphldf:hover, .p9NqC.kphldf:active { --gm-iconbutton-ink-color: var(--dt-error-action-stateful,rgb(179,20,18)); }

.p9NqC.kphldf:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.rNe0id { --mdc-ripple-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); --gm-iconbutton-ink-color: var(--dt-warning-action,rgb(60,64,67)); }

.p9NqC.rNe0id:focus, .p9NqC.rNe0id:hover, .p9NqC.rNe0id:active { --gm-iconbutton-ink-color: var(--dt-warning-action-stateful,rgb(32,33,36)); }

.p9NqC.rNe0id:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.sj692e { --mdc-ripple-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); --gm-iconbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); }

.p9NqC.sj692e:focus, .p9NqC.sj692e:hover, .p9NqC.sj692e:active { --gm-iconbutton-ink-color: var(--dt-primary-action-stateful,rgb(24,90,188)); }

.p9NqC.sj692e:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.IY5c4e { --mdc-ripple-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); --gm-iconbutton-ink-color: var(--dt-tertiary-action,rgb(19,115,51)); }

.p9NqC.IY5c4e:focus, .p9NqC.IY5c4e:hover, .p9NqC.IY5c4e:active { --gm-iconbutton-ink-color: var(--dt-tertiary-action-stateful,rgb(13,101,45)); }

.p9NqC.IY5c4e:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.qoCZef { --mdc-ripple-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); --gm-iconbutton-ink-color: var(--dt-neutral-action,rgb(60,64,67)); }

.p9NqC.qoCZef:focus, .p9NqC.qoCZef:hover, .p9NqC.qoCZef:active { --gm-iconbutton-ink-color: var(--dt-neutral-action-stateful,rgb(32,33,36)); }

.p9NqC.qoCZef:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.bustDd.sj692e, .p9NqC.bustDd.paynGb { --mdc-ripple-color: var(--dt-on-primary,#fff); --gm-iconbutton-ink-color: var(--dt-on-primary,#fff); }

.p9NqC.bustDd.sj692e:focus, .p9NqC.bustDd.sj692e:hover, .p9NqC.bustDd.sj692e:active, .p9NqC.bustDd.paynGb:focus, .p9NqC.bustDd.paynGb:hover, .p9NqC.bustDd.paynGb:active { --gm-iconbutton-ink-color: var(--dt-on-primary,#fff); }

.p9NqC.bustDd.sj692e:not(:disabled), .p9NqC.bustDd.paynGb:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.bustDd.IY5c4e { --mdc-ripple-color: var(--dt-on-tertiary,#fff); --gm-iconbutton-ink-color: var(--dt-on-tertiary,#fff); }

.p9NqC.bustDd.IY5c4e:focus, .p9NqC.bustDd.IY5c4e:hover, .p9NqC.bustDd.IY5c4e:active { --gm-iconbutton-ink-color: var(--dt-on-tertiary,#fff); }

.p9NqC.bustDd.IY5c4e:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.bustDd.qoCZef { --mdc-ripple-color: var(--dt-on-neutral,#fff); --gm-iconbutton-ink-color: var(--dt-on-neutral,#fff); }

.p9NqC.bustDd.qoCZef:focus, .p9NqC.bustDd.qoCZef:hover, .p9NqC.bustDd.qoCZef:active { --gm-iconbutton-ink-color: var(--dt-on-neutral,#fff); }

.p9NqC.bustDd.qoCZef:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.bustDd.kphldf { --mdc-ripple-color: var(--dt-on-error,#fff); --gm-iconbutton-ink-color: var(--dt-on-error,#fff); }

.p9NqC.bustDd.kphldf:focus, .p9NqC.bustDd.kphldf:hover, .p9NqC.bustDd.kphldf:active { --gm-iconbutton-ink-color: var(--dt-on-error,#fff); }

.p9NqC.bustDd.kphldf:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC.bustDd.rNe0id { --mdc-ripple-color: var(--dt-on-warning,rgb(32,33,36)); --gm-iconbutton-ink-color: var(--dt-on-warning,rgb(32,33,36)); }

.p9NqC.bustDd.rNe0id:focus, .p9NqC.bustDd.rNe0id:hover, .p9NqC.bustDd.rNe0id:active { --gm-iconbutton-ink-color: var(--dt-on-warning,rgb(32,33,36)); }

.p9NqC.bustDd.rNe0id:not(:disabled) { color: var(--gm-iconbutton-ink-color); }

.p9NqC:disabled { color: var(--dt-on-disabled,rgba(60,64,67,.38)); }

.usP4bb.kphldf { --gm-neutraltextbutton-ink-color: var(--dt-secondary-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-error-action-state-layer,rgb(197,34,31)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-error-action-stateful,rgb(179,20,18)); }

.usP4bb.rNe0id { --gm-neutraltextbutton-ink-color: var(--dt-secondary-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-warning-action-stateful,rgb(32,33,36)); }

.usP4bb.sj692e { --gm-neutraltextbutton-ink-color: var(--dt-secondary-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); }

.usP4bb.IY5c4e { --gm-neutraltextbutton-ink-color: var(--dt-secondary-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-tertiary-action-stateful,rgb(13,101,45)); }

.usP4bb.qoCZef { --gm-neutraltextbutton-ink-color: var(--dt-secondary-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-neutral-action-stateful,rgb(32,33,36)); }

.vhoiae .usP4bb.kphldf, .X9XeLb .usP4bb.kphldf, .cWKK1c .usP4bb.kphldf, .aJfoSc .usP4bb.kphldf, .TOb6Ze .usP4bb.kphldf { --gm-neutraltextbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-neutraltextbutton-state-color: var(--dt-error-action-state-layer,rgb(197,34,31)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-error-action-stateful,rgb(179,20,18)); }

.vhoiae .usP4bb.rNe0id, .X9XeLb .usP4bb.rNe0id, .cWKK1c .usP4bb.rNe0id, .aJfoSc .usP4bb.rNe0id, .TOb6Ze .usP4bb.rNe0id { --gm-neutraltextbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-neutraltextbutton-state-color: var(--dt-warning-action-state-layer,rgb(234,134,0)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-warning-action-stateful,rgb(32,33,36)); }

.vhoiae .usP4bb.sj692e, .X9XeLb .usP4bb.sj692e, .cWKK1c .usP4bb.sj692e, .aJfoSc .usP4bb.sj692e, .TOb6Ze .usP4bb.sj692e { --gm-neutraltextbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-neutraltextbutton-state-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); }

.vhoiae .usP4bb.IY5c4e, .X9XeLb .usP4bb.IY5c4e, .cWKK1c .usP4bb.IY5c4e, .aJfoSc .usP4bb.IY5c4e, .TOb6Ze .usP4bb.IY5c4e { --gm-neutraltextbutton-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-neutraltextbutton-state-color: var(--dt-tertiary-action-state-layer,rgb(19,115,51)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-tertiary-action-stateful,rgb(13,101,45)); }

.vhoiae .usP4bb.qoCZef, .X9XeLb .usP4bb.qoCZef, .cWKK1c .usP4bb.qoCZef, .aJfoSc .usP4bb.qoCZef, .TOb6Ze .usP4bb.qoCZef { --gm-neutraltextbutton-ink-color: var(--dt-neutral-action,rgb(60,64,67)); --gm-neutraltextbutton-state-color: var(--dt-neutral-action-state-layer,rgb(60,64,67)); --gm-neutraltextbutton-ink-color--stateful: var(--dt-neutral-action-stateful,rgb(32,33,36)); }

.vhoiae .xFWpbf.CZCFtc-bMElCd, .X9XeLb .xFWpbf.CZCFtc-bMElCd, .cWKK1c .xFWpbf.CZCFtc-bMElCd, .aJfoSc .xFWpbf.CZCFtc-bMElCd, .TOb6Ze .xFWpbf.CZCFtc-bMElCd { min-height: 2.5rem; }

.xFWpbf.CZCFtc-R6PoUb { height: 32px; margin-top: 0px; margin-bottom: 0px; }

.xFWpbf.CZCFtc-R6PoUb .VfPpkd-RLmnJb { height: 100%; }

.vhoiae .xFWpbf.CZCFtc-R6PoUb, .X9XeLb .xFWpbf.CZCFtc-R6PoUb, .cWKK1c .xFWpbf.CZCFtc-R6PoUb, .aJfoSc .xFWpbf.CZCFtc-R6PoUb, .TOb6Ze .xFWpbf.CZCFtc-R6PoUb { min-height: 2.25rem; }

.xFWpbf.CZCFtc-ibL1re { height: 28px; margin-top: 0px; margin-bottom: 0px; }

.xFWpbf.CZCFtc-ibL1re .VfPpkd-RLmnJb { height: 100%; }

.vhoiae .xFWpbf.CZCFtc-ibL1re, .X9XeLb .xFWpbf.CZCFtc-ibL1re, .cWKK1c .xFWpbf.CZCFtc-ibL1re, .aJfoSc .xFWpbf.CZCFtc-ibL1re, .TOb6Ze .xFWpbf.CZCFtc-ibL1re { min-height: 2rem; }

.xFWpbf.CZCFtc-c5RTEf { height: 24px; margin-top: 0px; margin-bottom: 0px; }

.xFWpbf.CZCFtc-c5RTEf .VfPpkd-RLmnJb { height: 100%; }

.vhoiae .xFWpbf.CZCFtc-c5RTEf, .X9XeLb .xFWpbf.CZCFtc-c5RTEf, .cWKK1c .xFWpbf.CZCFtc-c5RTEf, .aJfoSc .xFWpbf.CZCFtc-c5RTEf, .TOb6Ze .xFWpbf.CZCFtc-c5RTEf { min-height: 1.5rem; }

.vhoiae .p9NqC.CZCFtc-bMElCd, .X9XeLb .p9NqC.CZCFtc-bMElCd, .cWKK1c .p9NqC.CZCFtc-bMElCd, .aJfoSc .p9NqC.CZCFtc-bMElCd, .TOb6Ze .p9NqC.CZCFtc-bMElCd { min-height: 2.5rem; min-width: 2.5rem; }

.p9NqC.CZCFtc-R6PoUb { width: 44px; height: 44px; padding: 10px; }

.p9NqC.CZCFtc-R6PoUb .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 44px; max-width: 44px; }

.p9NqC.CZCFtc-R6PoUb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 40px; height: 40px; margin: 2px; }

.p9NqC.CZCFtc-R6PoUb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 40px; max-width: 40px; }

.p9NqC.CZCFtc-R6PoUb .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 44px; left: 50%; width: 44px; transform: translate(-50%, -50%); }

.vhoiae .p9NqC.CZCFtc-R6PoUb, .X9XeLb .p9NqC.CZCFtc-R6PoUb, .cWKK1c .p9NqC.CZCFtc-R6PoUb, .aJfoSc .p9NqC.CZCFtc-R6PoUb, .TOb6Ze .p9NqC.CZCFtc-R6PoUb { min-height: 2.25rem; min-width: 2.25rem; }

.p9NqC.CZCFtc-ibL1re { width: 40px; height: 40px; padding: 8px; }

.p9NqC.CZCFtc-ibL1re .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 40px; max-width: 40px; }

.p9NqC.CZCFtc-ibL1re.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 40px; height: 40px; margin: 0px; }

.p9NqC.CZCFtc-ibL1re.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 40px; max-width: 40px; }

.p9NqC.CZCFtc-ibL1re .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 40px; left: 50%; width: 40px; transform: translate(-50%, -50%); }

.vhoiae .p9NqC.CZCFtc-ibL1re, .X9XeLb .p9NqC.CZCFtc-ibL1re, .cWKK1c .p9NqC.CZCFtc-ibL1re, .aJfoSc .p9NqC.CZCFtc-ibL1re, .TOb6Ze .p9NqC.CZCFtc-ibL1re { min-height: 2rem; min-width: 2rem; }

.p9NqC.CZCFtc-c5RTEf { width: 36px; height: 36px; padding: 6px; }

.p9NqC.CZCFtc-c5RTEf .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 36px; max-width: 36px; }

.p9NqC.CZCFtc-c5RTEf.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 36px; height: 36px; margin: 0px; }

.p9NqC.CZCFtc-c5RTEf.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 36px; max-width: 36px; }

.p9NqC.CZCFtc-c5RTEf .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 36px; left: 50%; width: 36px; transform: translate(-50%, -50%); }

.vhoiae .p9NqC.CZCFtc-c5RTEf, .X9XeLb .p9NqC.CZCFtc-c5RTEf, .cWKK1c .p9NqC.CZCFtc-c5RTEf, .aJfoSc .p9NqC.CZCFtc-c5RTEf, .TOb6Ze .p9NqC.CZCFtc-c5RTEf { min-height: 1.5rem; min-width: 1.5rem; }

.p9NqC.CZCFtc-II5mzb { width: 32px; height: 32px; padding: 4px; }

.p9NqC.CZCFtc-II5mzb .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 32px; max-width: 32px; }

.p9NqC.CZCFtc-II5mzb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 32px; height: 32px; margin: 0px; }

.p9NqC.CZCFtc-II5mzb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 32px; max-width: 32px; }

.p9NqC.CZCFtc-II5mzb .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 32px; left: 50%; width: 32px; transform: translate(-50%, -50%); }

.p9NqC.CZCFtc-wNfPc { width: 28px; height: 28px; padding: 2px; }

.p9NqC.CZCFtc-wNfPc .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 28px; max-width: 28px; }

.p9NqC.CZCFtc-wNfPc.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc { width: 28px; height: 28px; margin: 0px; }

.p9NqC.CZCFtc-wNfPc.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec { max-height: 28px; max-width: 28px; }

.p9NqC.CZCFtc-wNfPc .VfPpkd-Bz112c-RLmnJb { position: absolute; top: 50%; height: 28px; left: 50%; width: 28px; transform: translate(-50%, -50%); }

.p9NqC.CZCFtc-wNfPc [viewbox] { height: 20px; padding: 2px; width: 20px; }

.cXSt5b:not(.JBW83d) { -webkit-box-align: center; align-items: center; display: flex; height: 18px; margin: 0px 8px 0px 0px; width: 18px; }

.cXSt5b.ZYNFl { margin: 0px 0px 0px 8px; }

.cXSt5b .mig17c { margin-left: -3px; }

html[dir="rtl"] .giSqbe { transform: scaleX(-1); }

.DU29of { position: relative; }

.DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo, .DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(66, 133, 244); }

@media screen and (forced-colors: active), (-ms-high-contrast:active) {
  .DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo, .DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(66, 133, 244); }

@media screen and (forced-colors: active), (-ms-high-contrast:active) {
  .DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(234, 67, 53); }

@media screen and (forced-colors: active), (-ms-high-contrast:active) {
  .DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(251, 188, 4); }

@media screen and (forced-colors: active), (-ms-high-contrast:active) {
  .DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: rgb(52, 168, 83); }

@media screen and (forced-colors: active), (-ms-high-contrast:active) {
  .DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G { stroke: canvastext; }
}

.DU29of .VfPpkd-JGcpL-Mr8B3-V67aGc { height: 100%; width: 100%; position: absolute; opacity: 0; overflow: hidden; z-index: -1; }

.AcBSlf { color: var(--dt-tertiary,rgb(24,128,56)); }

.f9rjnb, .uOObG { color: var(--dt-error,rgb(217,48,37)); }

.CUfc8e, .Ezbpyc { color: var(--dt-on-surface,rgb(60,64,67)); }

.OSbCNe { fill: var(--dt-primary,rgb(26,115,232)); }

.AeCFae, .L7BfGe { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.AeCFae { transform: rotate(0deg); }

.xapwh circle { fill: var(--dt-on-tertiary-container,rgb(60,64,67)); }

.xapwh path { fill: var(--dt-tertiary-container,rgb(230,244,234)); }

.rwb2Wb circle { fill: var(--dt-on-error-container,rgb(60,64,67)); }

.rwb2Wb path { fill: var(--dt-error-container,rgb(252,232,230)); }

.hotT5b circle { fill: transparent; }

.hotT5b path { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.k8ReU { fill: var(--dt-error,rgb(217,48,37)); }

.RAGhKc { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.uTs3jf { display: flex; justify-content: space-around; margin-top: 30%; width: 100%; }

.l5nOkf { fill: var(--dt-primary,rgb(26,115,232)); }

.GfKfSb { font-variant-numeric: tabular-nums; }

.UF1uUe { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.CBp5De { display: inline; }

.CBp5De .GfKfSb, .CBp5De .GfKfSb:not(:disabled) { border-radius: 80px; }

.WRrz1, .vxVgOe, .ujU03e { font-size: 14px; }

.WRrz1 { color: var(--dt-error,rgb(217,48,37)); fill: currentcolor; }

.vxVgOe { color: var(--dt-tertiary,rgb(24,128,56)); fill: currentcolor; }

.ujU03e { color: var(--dt-on-surface,rgb(60,64,67)); fill: currentcolor; }

.xocih { user-select: text; }

.d0RAsd { font: var(--dt-title-small-font,500 .875rem/1.25rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-small-spacing,.0178571429em); vertical-align: middle; }

.htwnvf .d0RAsd { text-decoration: line-through; }

.Gb84Ld { border-radius: var(--dt-corner-button,.25rem); margin-right: 8px; }

.lGln3c.eJxL0c.sZwqu { color: var(--dt-on-primary,#fff); background-color: rgb(26, 115, 232); }

.cYKmOb.eJxL0c.sZwqu:focus, .qEH5Fd.eJxL0c.sZwqu:focus, .cR63xd.eJxL0c.sZwqu:focus { background-color: rgb(27, 95, 185); }

.cYKmOb.eJxL0c.sZwqu::after, .qEH5Fd.eJxL0c.sZwqu::after, .cR63xd.eJxL0c.sZwqu::after { border-color: rgb(26, 115, 232); }

.cYKmOb.eJxL0c.sZwqu:hover, .qEH5Fd.eJxL0c.sZwqu:hover, .cR63xd.eJxL0c.sZwqu:hover { background-color: rgb(27, 102, 201); }

.cYKmOb.eJxL0c.sZwqu:active, .qEH5Fd.eJxL0c.sZwqu:active, .cR63xd.eJxL0c.sZwqu:active { background-color: rgb(27, 99, 193); }

.lGln3c.eJxL0c.pebthf { color: var(--dt-on-primary,#fff); background-color: rgb(217, 48, 37); }

.cYKmOb.eJxL0c.pebthf:focus, .qEH5Fd.eJxL0c.pebthf:focus, .cR63xd.eJxL0c.pebthf:focus { background-color: rgb(173, 44, 37); }

.cYKmOb.eJxL0c.pebthf::after, .qEH5Fd.eJxL0c.pebthf::after, .cR63xd.eJxL0c.pebthf::after { border-color: rgb(217, 48, 37); }

.cYKmOb.eJxL0c.pebthf:hover, .qEH5Fd.eJxL0c.pebthf:hover, .cR63xd.eJxL0c.pebthf:hover { background-color: rgb(187, 46, 37); }

.cYKmOb.eJxL0c.pebthf:active, .qEH5Fd.eJxL0c.pebthf:active, .cR63xd.eJxL0c.pebthf:active { background-color: rgb(180, 45, 37); }

.lGln3c.eJxL0c.scUZ3e { background-color: rgb(251, 188, 4); color: var(--dt-on-warning,rgb(32,33,36)); }

.cYKmOb.eJxL0c.scUZ3e:focus, .qEH5Fd.eJxL0c.scUZ3e:focus, .cR63xd.eJxL0c.scUZ3e:focus { background-color: rgb(198, 151, 12); }

.cYKmOb.eJxL0c.scUZ3e::after, .qEH5Fd.eJxL0c.scUZ3e::after, .cR63xd.eJxL0c.scUZ3e::after { border-color: rgb(251, 188, 4); }

.cYKmOb.eJxL0c.scUZ3e:hover, .qEH5Fd.eJxL0c.scUZ3e:hover, .cR63xd.eJxL0c.scUZ3e:hover { background-color: rgb(216, 163, 9); }

.cYKmOb.eJxL0c.scUZ3e:active, .qEH5Fd.eJxL0c.scUZ3e:active, .cR63xd.eJxL0c.scUZ3e:active { background-color: rgb(207, 157, 10); }

.lGln3c.eJxL0c.HQGKjb { color: var(--dt-on-primary,#fff); background-color: rgb(30, 142, 62); }

.cYKmOb.eJxL0c.HQGKjb:focus, .qEH5Fd.eJxL0c.HQGKjb:focus, .cR63xd.eJxL0c.HQGKjb:focus { background-color: rgb(30, 116, 56); }

.cYKmOb.eJxL0c.HQGKjb::after, .qEH5Fd.eJxL0c.HQGKjb::after, .cR63xd.eJxL0c.HQGKjb::after { border-color: rgb(30, 142, 62); }

.cYKmOb.eJxL0c.HQGKjb:hover, .qEH5Fd.eJxL0c.HQGKjb:hover, .cR63xd.eJxL0c.HQGKjb:hover { background-color: rgb(30, 125, 58); }

.cYKmOb.eJxL0c.HQGKjb:active, .qEH5Fd.eJxL0c.HQGKjb:active, .cR63xd.eJxL0c.HQGKjb:active { background-color: rgb(30, 120, 57); }

.lGln3c.eJxL0c.lQ3Lbf { color: var(--dt-on-primary,#fff); background-color: rgb(32, 33, 36); }

.cYKmOb.eJxL0c.lQ3Lbf:focus, .qEH5Fd.eJxL0c.lQ3Lbf:focus, .cR63xd.eJxL0c.lQ3Lbf:focus { background-color: rgb(86, 86, 89); }

.cYKmOb.eJxL0c.lQ3Lbf::after, .qEH5Fd.eJxL0c.lQ3Lbf::after, .cR63xd.eJxL0c.lQ3Lbf::after { border-color: rgb(32, 33, 36); }

.cYKmOb.eJxL0c.lQ3Lbf:hover, .qEH5Fd.eJxL0c.lQ3Lbf:hover, .cR63xd.eJxL0c.lQ3Lbf:hover { background-color: rgb(68, 69, 71); }

.cYKmOb.eJxL0c.lQ3Lbf:active, .qEH5Fd.eJxL0c.lQ3Lbf:active, .cR63xd.eJxL0c.lQ3Lbf:active { background-color: rgb(77, 77, 80); }

.lGln3c.VLrnY.sZwqu { color: rgb(24, 90, 188); background-color: rgb(232, 240, 254); }

.cYKmOb.VLrnY.sZwqu:focus, .qEH5Fd.VLrnY.sZwqu:focus, .cR63xd.VLrnY.sZwqu:focus { background-color: rgb(207, 222, 246); }

.cYKmOb.VLrnY.sZwqu::after, .qEH5Fd.VLrnY.sZwqu::after, .cR63xd.VLrnY.sZwqu::after { border-color: rgb(24, 90, 188); }

.cYKmOb.VLrnY.sZwqu:hover, .qEH5Fd.VLrnY.sZwqu:hover, .cR63xd.VLrnY.sZwqu:hover { background-color: rgb(224, 234, 251); }

.cYKmOb.VLrnY.sZwqu:active, .qEH5Fd.VLrnY.sZwqu:active, .cR63xd.VLrnY.sZwqu:active { background-color: rgb(211, 225, 247); }

.lGln3c.VLrnY.pebthf { color: rgb(179, 20, 18); background-color: rgb(252, 232, 230); }

.cYKmOb.VLrnY.pebthf:focus, .qEH5Fd.VLrnY.pebthf:focus, .cR63xd.VLrnY.pebthf:focus { background-color: rgb(243, 207, 205); }

.cYKmOb.VLrnY.pebthf::after, .qEH5Fd.VLrnY.pebthf::after, .cR63xd.VLrnY.pebthf::after { border-color: rgb(179, 20, 18); }

.cYKmOb.VLrnY.pebthf:hover, .qEH5Fd.VLrnY.pebthf:hover, .cR63xd.VLrnY.pebthf:hover { background-color: rgb(249, 224, 222); }

.cYKmOb.VLrnY.pebthf:active, .qEH5Fd.VLrnY.pebthf:active, .cR63xd.VLrnY.pebthf:active { background-color: rgb(245, 211, 209); }

.lGln3c.VLrnY.scUZ3e { color: rgb(32, 33, 36); background-color: rgb(254, 239, 195); }

.cYKmOb.VLrnY.scUZ3e:focus, .qEH5Fd.VLrnY.scUZ3e:focus, .cR63xd.VLrnY.scUZ3e:focus { background-color: rgb(227, 214, 176); }

.cYKmOb.VLrnY.scUZ3e::after, .qEH5Fd.VLrnY.scUZ3e::after, .cR63xd.VLrnY.scUZ3e::after { border-color: rgb(32, 33, 36); }

.cYKmOb.VLrnY.scUZ3e:hover, .qEH5Fd.VLrnY.scUZ3e:hover, .cR63xd.VLrnY.scUZ3e:hover { background-color: rgb(245, 231, 189); }

.cYKmOb.VLrnY.scUZ3e:active, .qEH5Fd.VLrnY.scUZ3e:active, .cR63xd.VLrnY.scUZ3e:active { background-color: rgb(232, 218, 179); }

.lGln3c.VLrnY.scUZ3e .daZhsc { color: rgb(227, 116, 0); }

.lGln3c.VLrnY.HQGKjb { color: rgb(19, 115, 51); background-color: rgb(230, 244, 234); }

.cYKmOb.VLrnY.HQGKjb:focus, .qEH5Fd.VLrnY.HQGKjb:focus, .cR63xd.VLrnY.HQGKjb:focus { background-color: rgb(205, 229, 212); }

.cYKmOb.VLrnY.HQGKjb::after, .qEH5Fd.VLrnY.HQGKjb::after, .cR63xd.VLrnY.HQGKjb::after { border-color: rgb(19, 115, 51); }

.cYKmOb.VLrnY.HQGKjb:hover, .qEH5Fd.VLrnY.HQGKjb:hover, .cR63xd.VLrnY.HQGKjb:hover { background-color: rgb(222, 239, 227); }

.cYKmOb.VLrnY.HQGKjb:active, .qEH5Fd.VLrnY.HQGKjb:active, .cR63xd.VLrnY.HQGKjb:active { background-color: rgb(209, 231, 216); }

.lGln3c.VLrnY.lQ3Lbf { color: rgb(32, 33, 36); background-color: rgb(241, 243, 244); }

.cYKmOb.VLrnY.lQ3Lbf:focus, .qEH5Fd.VLrnY.lQ3Lbf:focus, .cR63xd.VLrnY.lQ3Lbf:focus { background-color: rgb(216, 218, 219); }

.cYKmOb.VLrnY.lQ3Lbf::after, .qEH5Fd.VLrnY.lQ3Lbf::after, .cR63xd.VLrnY.lQ3Lbf::after { border-color: rgb(32, 33, 36); }

.cYKmOb.VLrnY.lQ3Lbf:hover, .qEH5Fd.VLrnY.lQ3Lbf:hover, .cR63xd.VLrnY.lQ3Lbf:hover { background-color: rgb(233, 235, 236); }

.cYKmOb.VLrnY.lQ3Lbf:active, .qEH5Fd.VLrnY.lQ3Lbf:active, .cR63xd.VLrnY.lQ3Lbf:active { background-color: rgb(220, 222, 223); }

.lGln3c.I5JVbf.sZwqu { border-color: rgb(26, 115, 232); color: rgb(24, 90, 188); background-color: transparent; }

.cYKmOb.I5JVbf.sZwqu:focus, .qEH5Fd.I5JVbf.sZwqu:focus, .cR63xd.I5JVbf.sZwqu:focus { background-color: rgba(24, 90, 188, 0.12); }

.cYKmOb.I5JVbf.sZwqu::after, .qEH5Fd.I5JVbf.sZwqu::after, .cR63xd.I5JVbf.sZwqu::after { border-color: rgb(26, 115, 232); }

.cYKmOb.I5JVbf.sZwqu:hover, .qEH5Fd.I5JVbf.sZwqu:hover, .cR63xd.I5JVbf.sZwqu:hover { background-color: rgba(24, 90, 188, 0.04); }

.cYKmOb.I5JVbf.sZwqu:active, .qEH5Fd.I5JVbf.sZwqu:active, .cR63xd.I5JVbf.sZwqu:active { background-color: rgba(24, 90, 188, 0.1); }

.lGln3c.I5JVbf.pebthf { border-color: rgb(217, 48, 37); color: rgb(179, 20, 18); background-color: transparent; }

.cYKmOb.I5JVbf.pebthf:focus, .qEH5Fd.I5JVbf.pebthf:focus, .cR63xd.I5JVbf.pebthf:focus { background-color: rgba(179, 20, 18, 0.12); }

.cYKmOb.I5JVbf.pebthf::after, .qEH5Fd.I5JVbf.pebthf::after, .cR63xd.I5JVbf.pebthf::after { border-color: rgb(217, 48, 37); }

.cYKmOb.I5JVbf.pebthf:hover, .qEH5Fd.I5JVbf.pebthf:hover, .cR63xd.I5JVbf.pebthf:hover { background-color: rgba(179, 20, 18, 0.04); }

.cYKmOb.I5JVbf.pebthf:active, .qEH5Fd.I5JVbf.pebthf:active, .cR63xd.I5JVbf.pebthf:active { background-color: rgba(179, 20, 18, 0.1); }

.lGln3c.I5JVbf.scUZ3e { border-color: rgb(234, 134, 0); color: rgb(32, 33, 36); background-color: transparent; }

.cYKmOb.I5JVbf.scUZ3e:focus, .qEH5Fd.I5JVbf.scUZ3e:focus, .cR63xd.I5JVbf.scUZ3e:focus { background-color: rgba(234, 134, 0, 0.12); }

.cYKmOb.I5JVbf.scUZ3e::after, .qEH5Fd.I5JVbf.scUZ3e::after, .cR63xd.I5JVbf.scUZ3e::after { border-color: rgb(234, 134, 0); }

.cYKmOb.I5JVbf.scUZ3e:hover, .qEH5Fd.I5JVbf.scUZ3e:hover, .cR63xd.I5JVbf.scUZ3e:hover { background-color: rgba(234, 134, 0, 0.04); }

.cYKmOb.I5JVbf.scUZ3e:active, .qEH5Fd.I5JVbf.scUZ3e:active, .cR63xd.I5JVbf.scUZ3e:active { background-color: rgba(234, 134, 0, 0.1); }

.lGln3c.I5JVbf.scUZ3e .daZhsc { color: rgb(234, 134, 0); }

.lGln3c.I5JVbf.HQGKjb { border-color: rgb(30, 142, 62); color: rgb(19, 115, 51); background-color: transparent; }

.cYKmOb.I5JVbf.HQGKjb:focus, .qEH5Fd.I5JVbf.HQGKjb:focus, .cR63xd.I5JVbf.HQGKjb:focus { background-color: rgba(19, 115, 51, 0.12); }

.cYKmOb.I5JVbf.HQGKjb::after, .qEH5Fd.I5JVbf.HQGKjb::after, .cR63xd.I5JVbf.HQGKjb::after { border-color: rgb(30, 142, 62); }

.cYKmOb.I5JVbf.HQGKjb:hover, .qEH5Fd.I5JVbf.HQGKjb:hover, .cR63xd.I5JVbf.HQGKjb:hover { background-color: rgba(19, 115, 51, 0.04); }

.cYKmOb.I5JVbf.HQGKjb:active, .qEH5Fd.I5JVbf.HQGKjb:active, .cR63xd.I5JVbf.HQGKjb:active { background-color: rgba(19, 115, 51, 0.1); }

.lGln3c.I5JVbf.lQ3Lbf { border-color: rgb(32, 33, 36); color: rgb(32, 33, 36); background-color: transparent; }

.cYKmOb.I5JVbf.lQ3Lbf:focus, .qEH5Fd.I5JVbf.lQ3Lbf:focus, .cR63xd.I5JVbf.lQ3Lbf:focus { background-color: rgba(32, 33, 36, 0.12); }

.cYKmOb.I5JVbf.lQ3Lbf::after, .qEH5Fd.I5JVbf.lQ3Lbf::after, .cR63xd.I5JVbf.lQ3Lbf::after { border-color: rgb(32, 33, 36); }

.cYKmOb.I5JVbf.lQ3Lbf:hover, .qEH5Fd.I5JVbf.lQ3Lbf:hover, .cR63xd.I5JVbf.lQ3Lbf:hover { background-color: rgba(32, 33, 36, 0.04); }

.cYKmOb.I5JVbf.lQ3Lbf:active, .qEH5Fd.I5JVbf.lQ3Lbf:active, .cR63xd.I5JVbf.lQ3Lbf:active { background-color: rgba(32, 33, 36, 0.1); }

.HTa8dc { background: none; border: none; color: inherit; font-family: inherit; font-size: inherit; margin: 0px; outline: none; padding: 0px; position: relative; }

.lGln3c { -webkit-box-align: center; align-items: center; border-radius: 0.25rem; box-sizing: border-box; display: inline-flex; max-width: 11.25rem; position: relative; vertical-align: middle; }

.lGln3c.w0hkKb { height: 1rem; }

.lGln3c.lSLCF { height: 1.25rem; }

.lGln3c > :not(:first-child) { padding-left: 0.125rem; }

.lGln3c > :first-child { border-bottom-left-radius: 0.25rem; border-top-left-radius: 0.25rem; padding-left: 0.25rem; }

.lGln3c > :not(:last-child) { padding-right: 0.125rem; }

.lGln3c > :last-child { border-bottom-right-radius: 0.25rem; border-top-right-radius: 0.25rem; padding-right: 0.25rem; }

.mLMBud { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-label-large-spacing,.0178571429em); box-sizing: border-box; font-size: 0.75rem; max-width: 100%; min-width: 0px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.cYKmOb { min-width: 0px; }

.cR63xd, .qEH5Fd, .cYKmOb { cursor: pointer; }

.cR63xd::after, .qEH5Fd::after, .cYKmOb::after { border-radius: 0.1875rem; border: 0.125rem solid rgb(26, 115, 232); inset: -0.1875rem; box-shadow: rgb(255, 255, 255) 0px 0px 0px 0.0625rem inset; content: ""; display: none; pointer-events: none; position: absolute; z-index: 1; }

.cR63xd:focus::after, .qEH5Fd:focus::after, .cYKmOb:focus::after { display: block; }

.cR63xd:focus:not(:focus-visible)::after, .qEH5Fd:focus:not(:focus-visible)::after, .cYKmOb:focus:not(:focus-visible)::after { display: none; }

.qEH5Fd, .cYKmOb { height: 100%; }

.cR63xd .mLMBud, .cYKmOb .mLMBud { text-decoration: underline; }

.cR63xd::after, .qEH5Fd:first-child::after, .cYKmOb:first-child::after { border-bottom-left-radius: 0.4375rem; border-top-left-radius: 0.4375rem; }

.cR63xd::after, .qEH5Fd:last-child::after, .cYKmOb:last-child::after { border-bottom-right-radius: 0.4375rem; border-top-right-radius: 0.4375rem; }

.hj61s, .qEH5Fd { -webkit-box-align: center; align-items: center; display: flex; }

.daZhsc.vKmmhc { fill: currentcolor; font-size: 1rem; height: 1rem; line-height: 1rem; width: 1rem; }

.daZhsc.vKmmhc [viewbox] { height: 1rem; width: 1rem; }

.lGln3c { border-color: transparent; }

.lGln3c::before { border-color: inherit; border-radius: 0.25rem; border-style: solid; border-width: 0.0625rem; box-sizing: border-box; content: ""; height: 100%; pointer-events: none; position: absolute; width: 100%; z-index: 1; }

c-wiz { contain: style; }

c-wiz > c-data { display: none; }

c-wiz.rETSD { contain: none; }

c-wiz.Ubi8Z { contain: layout style; }

.SN5W1d { box-sizing: border-box; color: var(--dt-on-surface-variant,rgb(95,99,104)); font-size: 1rem; margin-bottom: calc(1.9em - 1px); padding-bottom: 1px; position: relative; width: 100%; z-index: 0; }

.SN5W1d.FyWfTd { margin-bottom: 0px; padding-bottom: 0px; }

.SN5W1d.CDELXb { color: var(--dt-on-surface,rgb(60,64,67)); }

.SN5W1d.iPMcJc { color: var(--dt-primary-action,rgb(25,103,210)); }

.SN5W1d.Jj6Lae { color: var(--dt-error-action,rgb(197,34,31)); }

.mdf2C { -webkit-box-align: center; align-items: center; box-sizing: border-box; display: inline-flex; min-height: inherit; padding: 0px 0.75em; position: relative; width: 100%; }

.q300Cf { -webkit-box-flex: 1; flex: 1 1 auto; }

.BYnPEd { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-small-spacing,.025em); bottom: calc(-1.9em + 1px); box-sizing: border-box; color: var(--dt-on-surface-variant,rgb(95,99,104)); display: flex; fill: var(--dt-on-surface-variant,rgb(95,99,104)); font-size: 0.75em; height: 1.9em; left: 0px; line-height: 1.4em; max-width: 100%; padding: 0.35em 1.5em 0.1em; position: absolute; right: 0px; }

.BYnPEd.FyWfTd { display: none; }

.YXkYWb { -webkit-box-align: center; align-items: center; align-self: stretch; display: flex; -webkit-box-pack: start; justify-content: flex-start; position: relative; width: 100%; }

.LFY2Ee { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); align-self: stretch; display: flex; -webkit-box-flex: 1; flex: 1 1 auto; font-size: 0.875em; min-height: inherit; min-width: 0px; padding: 0px 0.125em 0px 0.25em; position: relative; width: 100%; }

.SUjDzd { box-sizing: border-box; cursor: text; font-size: 1.145em; max-width: 100%; user-select: none; z-index: 1; }

@media (forced-colors: active) {
  .SUjDzd { color: graytext; }
}

.hVDDMd { display: block; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.QipISb { display: flex; }

.o8tTsf { outline: none; overflow: hidden; text-overflow: ellipsis; }

.X2sj3b { padding-left: 0.25em; padding-right: 0.5em; }

.lIx1yc { padding-left: 0.25em; }

.X2sj3b, .lIx1yc { -webkit-box-align: center; align-items: center; align-self: flex-start; box-sizing: border-box; color: inherit; display: inline-flex; fill: currentcolor; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-pack: center; justify-content: center; }

.BYnPEd.Jj6Lae, .X2sj3b.Jj6Lae, .lIx1yc.Jj6Lae, .X2sj3b.Jj6Lae.Jj6Lae [viewbox], .lIx1yc.Jj6Lae.Jj6Lae [viewbox] { color: var(--dt-error-action,rgb(197,34,31)); fill: currentcolor; }

@media (forced-colors: active) {
  .X2sj3b, .lIx1yc { color: canvastext; }
}

.g1g2W { padding-top: 0.34375rem; }

.SN5W1d.EwXqJf { min-height: 3.5em; }

.SN5W1d.NWlIHc { min-height: 3.25em; }

.SN5W1d.nsKVp { min-height: 3em; }

.SN5W1d.GND07b { min-height: 2.7em; }

.SN5W1d.SjheHf { min-height: 2.5em; }

.SN5W1d.HHWuM { min-height: 2.25em; }

.SUjDzd.EwXqJf { height: 3.5em; }

.SUjDzd.NWlIHc { height: 3.25em; }

.SUjDzd.nsKVp { height: 3em; }

.SUjDzd.GND07b { height: 2.7em; }

.SUjDzd.SjheHf { height: 2.5em; }

.SUjDzd.HHWuM { height: 2.25em; }

.X2sj3b.EwXqJf, .lIx1yc.EwXqJf { height: 3.5em; }

.X2sj3b.NWlIHc, .lIx1yc.NWlIHc { height: 3.25em; }

.X2sj3b.nsKVp, .lIx1yc.nsKVp { height: 3em; }

.X2sj3b.GND07b, .lIx1yc.GND07b { height: 2.7em; }

.X2sj3b.SjheHf, .lIx1yc.SjheHf { height: 2.5em; }

.X2sj3b.HHWuM, .lIx1yc.HHWuM { height: 2.25em; }

.yid0mf { background: var(--dt-surface-variant,rgb(241,243,244)); border-bottom: 1px solid currentcolor; border-radius: var(--dt-corner-field-filled,.375rem .375rem 0 0); color: currentcolor; }

.yid0mf:not(.T3YfFf)::after { transition: transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.yid0mf:hover { background: var(--dt-surface-variant,rgb(241,243,244)); }

.yid0mf:hover::before { background: var(--dt-secondary-action-state-layer,rgb(60,64,67)); border-radius: var(--dt-corner-field-filled,.375rem .375rem 0 0); content: ""; height: 100%; left: 0px; opacity: 0.08; position: absolute; right: 0px; }

.yid0mf::after { border-bottom: 2px solid currentcolor; bottom: -1px; content: ""; height: 2px; left: 0px; position: absolute; right: 0px; transform: scaleX(0); z-index: 0; }

.yid0mf.Jj6Lae::after, .yid0mf.iPMcJc::after, .yid0mf.CDELXb::after { transform: scaleX(1); }

.yid0mf.Jj6Lae::after { border-color: var(--dt-error-action,rgb(197,34,31)); }

.yid0mf.iPMcJc { outline: transparent solid 1px; }

@media screen and (-ms-high-contrast:active) {
  .yid0mf { border-bottom-width: 2px; }
}

@media (forced-colors: active) {
  .yid0mf { border-bottom-color: buttontext; border-bottom-width: 1px; }
  .yid0mf::after { content: unset; transition: unset; }
  .yid0mf.iPMcJc, .yid0mf:hover { border-color: canvas; outline: none; }
  .yid0mf.iPMcJc::before, .yid0mf:hover::before { border-radius: inherit; border: 2px solid highlight; inset: 0px 0px -1px; content: ""; pointer-events: none; position: absolute; }
  .yid0mf.iPMcJc::after, .yid0mf:hover::after { border-radius: calc(var(--dt-corner-field-filled, .375rem .375rem 0 0) - 2px); border: 1px solid highlighttext; inset: 2px 2px 1px; content: ""; height: unset; pointer-events: none; position: absolute; transform: unset; z-index: unset; }
}

.DWM0ae { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-large-spacing,.00625em); -webkit-box-align: center; align-items: center; color: currentcolor; display: flex; font-size: 1.145em; left: 0.25em; pointer-events: none; position: absolute; top: 0px; transform: translateY(0px) scale(1); transform-origin: left top; }

.DWM0ae.iPMcJc, .DWM0ae.CDELXb { cursor: default; }

@media (forced-colors: active) {
  .DWM0ae { color: graytext; }
}

.xXpt7b.kM7Sgc.EwXqJf { padding-top: 1.35em; }

.xXpt7b.kM7Sgc.NWlIHc { padding-top: 1.3em; }

.xXpt7b.kM7Sgc.nsKVp { padding-top: 1.25em; }

.xXpt7b.kM7Sgc.GND07b { padding-top: 1.2em; }

.xXpt7b.kM7Sgc.SjheHf { padding-top: 1em; }

.DWM0ae:not(.T3YfFf) { transition: transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, color 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.DWM0ae.CDELXb, .DWM0ae.IbzNie, .DWM0ae.iPMcJc { transform: translateY(-10%) scale(0.75); }

.DWM0ae.VENvFd.iPMcJc { color: rgb(232, 113, 10); }

.xjBc3b { border: 1px solid var(--dt-outline,rgb(128,134,139)); border-radius: var(--dt-corner-field,.375rem); }

.xjBc3b::before { border: 1px solid transparent; border-radius: inherit; inset: -1px; content: ""; pointer-events: none; position: absolute; }

.xjBc3b:not(.T3YfFf)::before { transition: border 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.xjBc3b:hover::before { border-color: var(--dt-on-background,rgb(60,64,67)); }

.xjBc3b.ORw07d:hover::before { border-color: unset; }

.xjBc3b.iPMcJc::before, .xjBc3b.Jj6Lae::before { border: 2px solid currentcolor; }

.xjBc3b.Jj6Lae::before { border-color: var(--dt-error-action,rgb(197,34,31)); }

@media screen and (-ms-high-contrast:active) {
  .xjBc3b { border-width: 2px; }
}

@media (forced-colors: active) {
  .xjBc3b { border-color: buttontext; border-width: 1px; }
  .xjBc3b::before, .xjBc3b:hover::before { border-color: buttontext; transition: unset; }
  .xjBc3b.xjBc3b.xjBc3b::before { transition: unset; }
  .xjBc3b.iPMcJc, .xjBc3b:hover { border-color: canvas; outline: none; }
  .xjBc3b.iPMcJc::before, .xjBc3b:hover::before { border: 2px solid highlight; content: ""; }
  .xjBc3b.iPMcJc::after, .xjBc3b:hover::after { border-radius: calc(var(--dt-corner-field, .375rem) - 2px); border: 1px solid highlighttext; inset: 1px; content: ""; pointer-events: none; position: absolute; }
}

.iq7lKd { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-large-spacing,.00625em); -webkit-box-align: center; align-items: center; box-sizing: border-box; bottom: 0px; color: currentcolor; display: flex; font-size: 1.145em; max-width: 100%; position: absolute; top: 0px; transform: translateX(-0.35em) scale(1); transform-origin: left top; }

.iq7lKd.iPMcJc, .iq7lKd.CDELXb { cursor: default; }

@media (forced-colors: active) {
  .iq7lKd { color: graytext; }
}

.iq7lKd.Jj6Lae.iPMcJc { color: var(--dt-error-action,rgb(197,34,31)); }

.tknroe { box-sizing: border-box; overflow: hidden; padding: 0px 0.25em; }

.iq7lKd:not(.T3YfFf) { transition: transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, max-width 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, color 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.iq7lKd.CDELXb, .iq7lKd.IbzNie, .iq7lKd.iPMcJc { transform: translateY(-36%) scale(0.75); max-width: 133%; }

.CeSLIf { background: linear-gradient(180deg,var(--dt-background,#fff) 0,var(--dt-background,#fff) 70%,transparent 70%,transparent 100%); padding: 0px 0.25em; }

@media (forced-colors: active) {
  .CeSLIf { background: none; }
}

.RE1Byf { background: var(--dt-surface-variant,rgb(241,243,244)); border: 1px solid transparent; border-radius: var(--dt-corner-field-search,.5rem); box-shadow: none; }

.vhoiae .RE1Byf, .X9XeLb .RE1Byf, .cWKK1c .RE1Byf, .aJfoSc .RE1Byf, .TOb6Ze .RE1Byf { background: var(--dt-surface3,#fff); }

.RE1Byf:hover { border-color: rgb(232, 234, 237); }

.RE1Byf.iPMcJc { background: var(--dt-surface1,#fff); box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.vhoiae .RE1Byf.iPMcJc, .X9XeLb .RE1Byf.iPMcJc, .cWKK1c .RE1Byf.iPMcJc, .aJfoSc .RE1Byf.iPMcJc, .TOb6Ze .RE1Byf.iPMcJc { background: var(--dt-surface,#fff); }

.RE1Byf.Jj6Lae { color: var(--dt-error-action,rgb(197,34,31)); }

@media screen and (-ms-high-contrast:active) {
  .RE1Byf { border: solid 2px var(--dt-outline,rgb(128,134,139)); }
  .RE1Byf:hover { border-color: rgb(95, 99, 104); }
  .RE1Byf.iPMcJc { border-color: var(--dt-primary-action,rgb(25,103,210)); }
}

@media (forced-colors: active) {
  .RE1Byf, .RE1Byf:hover { border-color: buttontext; border-width: 1px; }
  .RE1Byf.iPMcJc, .RE1Byf:hover { border-color: canvas; outline: none; }
  .RE1Byf.iPMcJc::before, .RE1Byf:hover::before { border-radius: inherit; border: 2px solid highlight; inset: -1px; content: ""; pointer-events: none; position: absolute; }
  .RE1Byf.iPMcJc::after, .RE1Byf:hover::after { border-radius: calc(var(--dt-corner-field-search, .5rem) - 2px); border: 1px solid highlighttext; inset: 1px; content: ""; pointer-events: none; position: absolute; }
}

.rj3NAb { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-body-large-spacing,.00625em); -webkit-box-align: center; align-items: center; bottom: 0px; color: var(--dt-on-surface-variant,rgb(95,99,104)); display: flex; font-size: 1.145em; left: 0.25ch; margin: 0px 0.15em; position: absolute; top: 0px; }

@media (forced-colors: active) {
  .rj3NAb { color: graytext; }
}

.rj3NAb.Jj6Lae { color: var(--dt-error-action,rgb(197,34,31)); }

.rj3NAb.CDELXb, .rj3NAb.IbzNie { display: none; }

.LUNIy { background: transparent; border: none; box-shadow: none; box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); display: inline-block; font-family: Roboto, Arial, sans-serif; font-size: 1em; margin: 0px; min-height: 1.75em; padding: 0.25em 0px; width: 100%; }

.LUNIy, .LUNIy:focus, .LUNIy:active { outline: none; }

.LUNIy.q4tg { outline: none; resize: none; overflow: hidden auto; }

.LUNIy.q4tg::-webkit-scrollbar { display: none; }

@-webkit-keyframes quantumWizBoxInkSpread { 
  0% { transform: translate(-50%, -50%) scale(0.2); }
  100% { transform: translate(-50%, -50%) scale(2.2); }
}

@keyframes quantumWizBoxInkSpread { 
  0% { transform: translate(-50%, -50%) scale(0.2); }
  100% { transform: translate(-50%, -50%) scale(2.2); }
}

@-webkit-keyframes quantumWizIconFocusPulse { 
  0% { transform: translate(-50%, -50%) scale(1.5); opacity: 0; }
  100% { transform: translate(-50%, -50%) scale(2); opacity: 1; }
}

@keyframes quantumWizIconFocusPulse { 
  0% { transform: translate(-50%, -50%) scale(1.5); opacity: 0; }
  100% { transform: translate(-50%, -50%) scale(2); opacity: 1; }
}

@-webkit-keyframes quantumWizRadialInkSpread { 
  0% { transform: scale(1.5); opacity: 0; }
  100% { transform: scale(2.5); opacity: 1; }
}

@keyframes quantumWizRadialInkSpread { 
  0% { transform: scale(1.5); opacity: 0; }
  100% { transform: scale(2.5); opacity: 1; }
}

@-webkit-keyframes quantumWizRadialInkFocusPulse { 
  0% { transform: scale(2); opacity: 0; }
  100% { transform: scale(2.5); opacity: 1; }
}

@keyframes quantumWizRadialInkFocusPulse { 
  0% { transform: scale(2); opacity: 0; }
  100% { transform: scale(2.5); opacity: 1; }
}

.OTFkff { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); height: 1.75rem; min-height: 40px; padding: 0.625rem 0px; outline: none; overflow: hidden; white-space: pre-wrap; width: 100%; overflow-wrap: break-word; }

.DpejEd { transition: opacity 0.2s ease-in-out 0s; opacity: 0; }

.DpejEd.aPfFOd { opacity: 1; }

.W6Pykc { margin: 0px -6px; }

.WyLv6c { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; }

.XQGDUc { display: flex; }

.ElDLFb { -webkit-box-align: center; align-items: center; display: flex; }

.ElDLFb.syTahf { width: auto; }

.cqt6tc { background: var(--dt-inverse-surface,rgb(32,33,36)); inset: 0px; display: none; opacity: 0.5; position: absolute; z-index: 1000; }

.XQGDUc[aria-expanded="true"] .cqt6tc { display: block; }

.XQGDUc .wr0Q1d.wr0Q1d { place-content: center flex-start; border-radius: var(--dt-corner-button,.25rem); box-sizing: border-box; -webkit-box-pack: start; overflow: hidden; padding: 6px 45px 6px 8px; }

.XQGDUc .wr0Q1d.syTahf { padding: 6px 14px 6px 8px; width: auto; }

.XQGDUc.L2G7g .wr0Q1d { border-radius: 16px; height: 32px; }

.XQGDUc.L2G7g .wr0Q1d.syTahf { display: none; }

.NqtXkd { align-self: center; fill: var(--dt-primary-action,rgb(25,103,210)); height: 18px; margin-right: 8px; width: 18px; }

.jfV46c { fill: var(--dt-primary-action,rgb(25,103,210)); }

.JQNYBe { -webkit-box-align: center; align-items: center; border-top: solid 1px var(--dt-outline-variant,rgb(218,220,224)); -webkit-box-pack: center; justify-content: center; padding: 6px 0px; }

.sQFJD { display: flex; }

.s7kctf, .SfRhr { align-self: center; display: flex; }

.eQcqZd { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.vG8rmc { color: var(--dt-on-surface-variant,rgb(95,99,104)); margin: 0px 18px 0px 14px; width: 100%; }

.Ot6Nnc { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 6px 6px 6px 0px; }

.XFWqvb { align-self: center; position: relative; right: 45px; }

.hDzJ7b { width: 250px; }

.Nh8zLd { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.wr0Q1d [jsname="label_"] { position: relative; top: 1px; }

.y0vmdf { -webkit-box-align: center; align-items: center; inset: 0px; display: flex; -webkit-box-pack: center; justify-content: center; position: absolute; z-index: 2000; }

.y0vmdf:not(.BXXR1b) { display: none; }

.R8blcc { background-color: rgba(0, 0, 0, 0.5); position: absolute; height: 100%; width: 100%; z-index: 1; }

.ZNusbb { background-color: var(--dt-surface3,#fff); border-radius: 8px; box-shadow: rgba(0, 0, 0, 0.2) 0px 1px 3px; width: 204px; padding: 25px; z-index: 2; }

.f1vfGd { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,.00625em); color: var(--dt-on-surface,rgb(60,64,67)); display: block; padding-bottom: 12px; }

.CflXCe { font: var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-large-spacing,.00625em); color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.F0AQmf.eLNT1d { display: none; }

.cNoHqf { width: 100%; }

.cNoHqf .snByac { z-index: 1; }

.cNoHqf .snByac .CeSLIf { background: linear-gradient(180deg,var(--dt-surface3,#fff) 0,var(--dt-surface3,#fff) 70%,transparent 70%,transparent 100%); }

.i1aqqc { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: end; justify-content: flex-end; padding-top: 18px; }

.YXvFRd { margin-right: 10px; }

.SNsaHc { fill: var(--dt-tertiary-icon,#fff); }

.AB2z5e { white-space: nowrap; }

.wichcb { appearance: none; -webkit-box-align: center; align-items: center; background: transparent; border: none; display: inline-flex; color: inherit; font-style: inherit; font-variant: inherit; font-weight: inherit; font-stretch: inherit; font-size: inherit; font-family: inherit; font-optical-sizing: inherit; font-kerning: inherit; font-feature-settings: inherit; font-variation-settings: inherit; -webkit-box-pack: center; justify-content: center; line-height: normal; margin: 0px; overflow: visible; padding: 0px; text-align: inherit; width: auto; }

.yQJ3f { box-sizing: border-box; border-radius: inherit; max-height: 100%; max-width: 100%; }

.igenxd { border-radius: inherit; display: inline-block; }

.EHUFff { -webkit-box-align: center; place-items: center start; box-sizing: border-box; display: grid; grid-template-columns: 1fr auto auto; padding: 0px 1.25rem 0px 0.5rem; height: 3.5rem; }

.zPuWle { display: none; }

.wQArwd { display: block; max-width: 100%; width: 100%; }

.CJiroe { display: grid; grid-template-columns: repeat(7, 1fr); height: 40px; }

.CJiroe.hncTuf { clip-path: inset(50%); clip: rect(1px, 1px, 1px, 1px); height: 1px; margin: -1px; opacity: 0; overflow: hidden; padding: 0px; position: absolute; width: 1px; }

.KtZAl { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); -webkit-box-align: center; align-items: center; box-sizing: border-box; display: flex; height: 40px; -webkit-box-pack: center; justify-content: center; width: 40px; }

.RwDu8c { background-color: var(--dt-surface,#fff); border-radius: inherit; color: var(--dt-on-surface,rgb(60,64,67)); position: relative; width: 296px; }

.RwDu8c > [role="listbox"] { outline: none; }

.GBsejc { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-weight: ; font-stretch: ; font-size: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-title-small-spacing,.0178571429em); border-radius: var(--dt-corner-button,.25rem); color: var(--dt-on-surface,rgb(60,64,67)); text-align: center; cursor: pointer; height: 1.75rem; line-height: 1.75rem; padding: 0px 1.25rem 0px 1rem; position: relative; }

.GBsejc::after { border-color: var(--dt-on-surface,rgb(60,64,67)) transparent; border-style: solid; border-width: 5px 4px 0px; bottom: 0px; content: " "; height: 4px; position: absolute; right: 6px; top: 12px; }

.tn62od { text-align: right; }

.Tx3nse { margin: 1px; }

.ZNYEy { color: var(--dt-on-surface,rgb(60,64,67)); }

.XjokOb { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); -webkit-box-align: center; align-items: center; box-sizing: border-box; border-radius: 50%; color: var(--dt-on-surface,rgb(60,64,67)); cursor: pointer; display: flex; -webkit-box-pack: center; justify-content: center; height: 100%; min-width: 100%; outline: none; padding: 0px; position: relative; text-align: center; vertical-align: middle; width: 100%; }

.XjokOb:focus { outline: none; }

.XjokOb.KKjvXb { background-color: var(--dt-primary,rgb(26,115,232)); color: var(--dt-on-primary,#fff); }

.XjokOb.RDPZE { color: var(--dt-on-disabled,rgba(60,64,67,.38)); cursor: default; }

.XjokOb.KKjvXb:not(:empty) { background: var(--dt-primary-action,rgb(25,103,210)); }

.XjokOb.KKjvXb:not(:empty)::before { border-radius: 50%; inset: 0px; content: ""; position: absolute; }

.XjokOb.KKjvXb:not(:empty)::before { border: 2px solid transparent; }

.DAx1Cc { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; max-height: 250px; overflow: hidden auto; }

.XvN0je { cursor: pointer; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; flex-shrink: 0; height: 40px; -webkit-box-pack: center; justify-content: center; text-align: center; width: 286px; }

.XvN0je[aria-disabled="true"] { color: var(--dt-on-disabled,rgba(60,64,67,.38)); }

@media screen and (forced-colors: active) {
  .XvN0je[aria-disabled="true"] { color: graytext; }
}

.XvN0je[aria-selected="true"] { font-size: 150%; }

.XvN0je.TrJ0Tc { color: var(--dt-primary-action,rgb(25,103,210)); font-size: 150%; }

.e431ed { cursor: pointer; }

.l8ICnb { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); display: block; outline: none; padding: 8px; }

.l8ICnb:focus { outline: none; }

.AAAnue { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.Ss7qXc { outline: none; position: relative; }

.Ss7qXc:focus { outline: none; }

.WNpj6b, .cUCuw { border-radius: inherit; box-sizing: border-box; color: currentcolor; display: none; font-style: normal; inset: 0px; position: absolute; pointer-events: none; }

.WNpj6b { border-radius: 0.375rem; border: .125rem solid var(--dt-primary-action-stateful,rgb(24,90,188)); z-index: 1; }

.WNpj6b::after { border-radius: 0.4375rem; border: .125rem solid var(--dt-primary-container,rgb(232,240,254)); content: ""; pointer-events: none; position: absolute; }

.WNpj6b.i1jHKe { inset: -0.25rem; }

.WNpj6b.i1jHKe::after { inset: -0.25rem; }

.WNpj6b.o1CAae { border-radius: inherit; inset: -0.25rem; }

.WNpj6b.o1CAae::after { border-radius: inherit; inset: -0.25rem; }

.WNpj6b.DMO9bd { inset: 0px; }

.WNpj6b.DMO9bd::after { inset: 0px; }

.WNpj6b.LwVLic { border-radius: inherit; inset: 0px; }

.WNpj6b.LwVLic::after { border-radius: inherit; inset: 0px; }

.cUCuw { background-color: currentcolor; z-index: 0; }

.Ss7qXc.Iryyw .cUCuw { z-index: -1; }

.Ss7qXc:hover .vA3Shd, .Ss7qXc.Iryyw :hover ~ .vA3Shd, .Ss7qXc.pBhGie .vA3Shd { opacity: 0.08; }

.Ss7qXc:active .upeNge, .Ss7qXc.Iryyw :active ~ .upeNge, .Ss7qXc.qs41qe .upeNge { opacity: 0.12; }

.Ss7qXc:focus .QmyJdb, .Ss7qXc.Iryyw :focus ~ .QmyJdb, .Ss7qXc.u3bW4e .QmyJdb { opacity: 0.12; }

.Ss7qXc[aria-grabbed="true"] .KuOzJf, .Ss7qXc.Iryyw [aria-grabbed="true"] ~ .KuOzJf, .Ss7qXc.MILgc .KuOzJf { opacity: 0.16; }

.Ss7qXc:active .upeNge, .Ss7qXc.qs41qe .upeNge, .Ss7qXc:focus .QmyJdb, .Ss7qXc.u3bW4e .QmyJdb, .Ss7qXc:focus-visible .WNpj6b, .Ss7qXc.GrxScd .WNpj6b, .Ss7qXc:hover .vA3Shd, .Ss7qXc.pBhGie .vA3Shd, .Ss7qXc.MILgc .KuOzJf, .Ss7qXc[aria-grabbed="true"] .KuOzJf { display: block; }

.Ss7qXc.Iryyw :focus-visible ~ .WNpj6b, .Ss7qXc.Iryyw :active ~ .upeNge, .Ss7qXc.Iryyw :focus ~ .QmyJdb, .Ss7qXc.Iryyw :hover ~ .vA3Shd, .Ss7qXc.Iryyw [aria-grabbed="true"] ~ .KuOzJf { display: block; }

.Ss7qXc:active .Ss7qXc:not(:active) .upeNge, .Ss7qXc.qs41qe .Ss7qXc:not(.qs41qe) .upeNge, .Ss7qXc:focus .Ss7qXc:not(:focus) .QmyJdb, .Ss7qXc.u3bW4e .Ss7qXc:not(.u3bW4e) .QmyJdb, .Ss7qXc:focus-visible .Ss7qXc:not(:focus-visible) .WNpj6b, .Ss7qXc.GrxScd .Ss7qXc:not(.GrxScd) .WNpj6b, .Ss7qXc:hover .Ss7qXc:not(:hover) .vA3Shd, .Ss7qXc.pBhGie .Ss7qXc:not(.pBhGie) .vA3Shd, .Ss7qXc.MILgc .Ss7qXc:not(.MILgc) .KuOzJf, .Ss7qXc[aria-grabbed="true"] .Ss7qXc[aria-grabbed="undefined"] .KuOzJf, .Ss7qXc[aria-grabbed="true"] .Ss7qXc[aria-grabbed="false"] .KuOzJf { display: none; }

.zAfnEf { background: var(--dt-surface,#fff); border-radius: var(--dt-corner-dialog-anchored,.5rem); box-shadow: var(--dt-surface3-shadow,0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15)); display: block; padding: 0px; position: absolute; width: 18.5rem; z-index: 2000; }

@media (forced-colors: active) {
  .zAfnEf { border: 1px solid canvastext; }
}

.zAfnEf.zmK2he { position: fixed; }

.zAfnEf:not(.eO2Zfd), .zAfnEf.BIIBbc { display: none; }

.M4Vw0b { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 1rem 1.5rem; }

.M4Vw0b:not(.eO2Zfd) { display: none; }

.oQSg1c { font: var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-large-spacing,0); color: var(--dt-on-surface,rgb(60,64,67)); padding: 1.5rem 1.5rem 0.5rem; }

.DuCDAf { inset: 0px; position: fixed; z-index: -1; }

.lvPJU { display: none; }

.HdS2Fc { background: transparent; border: 0px; color: inherit; margin: 0px; padding: 0px; vertical-align: baseline; }

.xz1uh { font-weight: 700; }

.C9D8j { list-style: none; margin: 0px; max-height: 100%; max-width: 100%; outline: none; padding: 0px; }

.C9D8j[aria-orientation="horizontal"] { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; }

.ia8caf { position: relative; }

.E4TL5c { position: absolute; left: 100%; top: 0px; }

.E4TL5c.eLNT1d { visibility: hidden; }

.E4TL5c.JGA0ke { left: auto; right: 100%; }

.ia8caf[aria-expanded="false"] .E4TL5c { pointer-events: none; opacity: 0; }

.eohZq { box-sizing: border-box; visibility: visible; max-height: 100%; max-width: 100%; z-index: 0; }

.gVl2db { background-color: var(--dt-surface3,#fff); border-radius: 8px; box-sizing: border-box; list-style: none; margin: 0px; max-width: 100%; min-width: 12rem; padding: 0.5rem 0px; position: relative; transform-origin: left top; z-index: 2300; }

.gVl2db:not(.AZSdVb) { max-height: 20rem; overflow-y: auto; }

.gVl2db:not(:empty) { box-shadow: var(--dt-surface2-shadow,0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)); }

.vhoiae .gVl2db { background: var(--dt-background,#fff); }

:not(.eLNT1d) > .gVl2db { animation: 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running menu-keyframes-zoom; }

[hidden] .eohZq { display: none; }

.Zw2DU { top: -0.5rem; }

.dT7Zpe { border-top: 1px solid var(--dt-outline,rgb(128,134,139)); height: 0px; margin: 0.375rem 0px; }

.b9OJXe { font: var(--dt-label-small-font,500 .6875rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-small-spacing,.0727272727em); text-transform: var(--dt-label-small-transform,uppercase); color: var(--dt-on-surface-variant,rgb(95,99,104)); padding: 0.75rem 1rem 0.5rem; }

.zycvZb, .tJCjXc { list-style: none; margin: 0px; padding: 0px; }

.WP8l3b { place-content: center; -webkit-box-align: center; align-items: center; box-sizing: border-box; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-pack: center; min-width: 3.25rem; }

.WP8l3b.JU2QSe { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.WP8l3b.JU2QSe.s4Oi9c { height: 1.25rem; padding: 0px 1rem; width: 1.25rem; }

.ZzDyt { -webkit-box-align: center; align-items: center; box-sizing: border-box; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-pack: end; justify-content: flex-end; margin: 0px 1rem; }

.rDy0g { text-transform: uppercase; }

.Wp3BKe { box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); font-size: 0.875rem; line-height: 1.25rem; list-style-image: none; outline: none; padding: 0px; position: relative; }

.Wp3BKe::before { inset: 0px; content: ""; position: absolute; }

.Wp3BKe:hover::before, .Wp3BKe:active::before { background: var(--dt-surface-variant,rgb(241,243,244)); }

.Wp3BKe:focus::before, .Wp3BKe.qs41qe::before, .Wp3BKe[aria-expanded="true"]::before { background: var(--dt-on-surface,rgb(60,64,67)); opacity: 0.12; }

.Wp3BKe[aria-selected="true"], .Wp3BKe[aria-checked="true"] { background: var(--dt-primary-container,rgb(232,240,254)); }

.Wp3BKe[aria-disabled], .Wp3BKe[disabled] { opacity: 0.38; }

.vUBIke { -webkit-box-align: center; align-items: center; background-color: transparent; box-sizing: border-box; display: flex; -webkit-box-pack: start; justify-content: flex-start; flex-wrap: nowrap; min-height: 22px; padding: 0.25rem 1rem; pointer-events: none; position: relative; z-index: 0; }

.vUBIke.glq6wf { padding-left: 0px; }

.vUBIke.mxtwQe { padding-right: 0px; }

.vUBIke.ncMAWe { min-height: 2.5rem; }

.vUBIke.ncMAWe.STFd6 { min-height: 3.75rem; }

.vUBIke.s4Oi9c { min-height: 2rem; }

.vUBIke.s4Oi9c.STFd6 { min-height: 3.25rem; }

.nYEsj { display: flex; -webkit-box-pack: center; justify-content: center; line-height: 0; overflow: hidden; }

.HWU5k { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; box-sizing: border-box; display: block; -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; letter-spacing: 0.2px; pointer-events: none; text-overflow: ellipsis; transform-style: preserve-3d; white-space: nowrap; }

.HWU5k.evOMld { text-overflow: clip; white-space: normal; word-break: break-word; }

.szjM5b { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); box-sizing: border-box; color: var(--dt-on-surface-variant,rgb(95,99,104)); display: block; overflow: hidden; text-decoration: inherit; text-overflow: ellipsis; text-transform: inherit; transform-style: preserve-3d; white-space: nowrap; }

.szjM5b.evOMld { text-overflow: clip; white-space: normal; word-break: break-word; }

@media (forced-colors: active) {
  .Wp3BKe[aria-disabled] .HWU5k, .Wp3BKe[disabled] .HWU5k, .Wp3BKe[aria-disabled] .szjM5b, .Wp3BKe[disabled] .szjM5b { color: graytext; }
}

@media (forced-colors: active) {
  .szjM5b.qs41qe, .HWU5k.qs41qe { color: highlighttext; }
}

.BWglse { display: block; height: 0px; overflow: hidden; width: 0px; }

.zoqPuc { color: var(--dt-primary,rgb(26,115,232)); }

.ZXFLTe { color: var(--dt-on-surface-variant,rgb(95,99,104)); height: 1.25rem; width: 1.25rem; }

.JhTOge { color: inherit; text-decoration: none; }

.JhTOge:focus { outline: none; }

@-webkit-keyframes menu-keyframes-zoom { 
  0% { opacity: 0; transform: scale(0.9); }
  30% { opacity: 1; }
  100% { opacity: 1; transform: none; }
}

@keyframes menu-keyframes-zoom { 
  0% { opacity: 0; transform: scale(0.9); }
  30% { opacity: 1; }
  100% { opacity: 1; transform: none; }
}

.FDSlxb.vf9sSe { border-radius: inherit; inset: 0px; display: block; pointer-events: auto; position: absolute; user-select: none; }

.KUcxMe .snByac { cursor: default; }

.Vf3OKe { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); background: none; border: none; color: var(--dt-on-surface,rgb(60,64,67)); min-height: 1.75em; outline: none; overflow: hidden; padding: 0px; text-align: left; text-overflow: ellipsis; white-space: nowrap; width: 100%; }

.Vf3OKe[aria-disabled="true"] { color: var(--dt-on-surface-secondary,rgb(95,99,104)); }

.Vf3OKe:focus { outline: none; }

@media (forced-colors: active) {
  .Vf3OKe, .Vf3OKe[aria-disabled="true"] { background-color: canvas; color: fieldtext; }
}

.i1wuu { vertical-align: middle; }

.f8KRkf { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,.0178571429em); }

.tqPe5c { color: var(--dt-primary,rgb(26,115,232)); }

.DPvwYc { font-family: "Material Icons Extended"; font-weight: normal; font-style: normal; font-size: 24px; line-height: 1; letter-spacing: normal; text-rendering: optimizelegibility; text-transform: none; display: inline-block; overflow-wrap: normal; direction: ltr; font-feature-settings: "liga"; -webkit-font-smoothing: antialiased; }

html[dir="rtl"] .sm8sCf { transform: scaleX(-1); }

.JPdR6b { transform: translateZ(0px); transition: max-width 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, max-height 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, opacity 0.1s linear 0s; background: rgb(255, 255, 255); border: 0px; border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; box-sizing: border-box; max-height: 100%; max-width: 100%; opacity: 1; outline: transparent solid 1px; z-index: 2000; }

.XvhY1d { overflow: hidden auto; }

.JAPqpe { float: left; padding: 16px 0px; }

.JPdR6b.qjTEB { transition: left 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, max-width 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, max-height 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, opacity 0.05s linear 0s, top 0.2s cubic-bezier(0, 0, 0.2, 1) 0s; }

.JPdR6b.jVwmLb { max-height: 56px; opacity: 0; }

.JPdR6b.CAwICe { overflow: hidden; }

.JPdR6b.oXxKqf { transition: none 0s ease 0s; }

.z80M1 { color: rgb(34, 34, 34); cursor: pointer; display: block; outline: none; overflow: hidden; padding: 0px 24px; position: relative; }

.uyYuVb { display: flex; font-size: 14px; font-weight: 400; line-height: 40px; height: 40px; position: relative; white-space: nowrap; }

.jO7h3c { -webkit-box-flex: 1; flex-grow: 1; min-width: 0px; }

.JPdR6b.e5Emjc .z80M1 { padding-left: 64px; }

.JPdR6b.CblTmf .z80M1 { padding-right: 48px; }

.PCdOIb { display: flex; flex-direction: column; justify-content: center; background-repeat: no-repeat; height: 40px; left: 24px; opacity: 0.54; position: absolute; }

.z80M1.RDPZE .PCdOIb { opacity: 0.26; }

.z80M1.FwR7Pc { outline: transparent solid 1px; background-color: rgb(238, 238, 238); }

.z80M1.RDPZE { color: rgb(184, 184, 184); cursor: default; }

.z80M1.N2RpBe::before { transform: rotate(45deg); transform-origin: left center; content: " "; display: block; border-right: 2px solid rgb(34, 34, 34); border-bottom: 2px solid rgb(34, 34, 34); height: 16px; left: 24px; opacity: 0.54; position: absolute; top: 13%; width: 7px; z-index: 0; }

.JPdR6b.CblTmf .z80M1.N2RpBe::before { left: auto; right: 16px; }

.z80M1.RDPZE::before { border-color: rgb(184, 184, 184); opacity: 1; }

.aBBjbd { pointer-events: none; position: absolute; }

.z80M1.qs41qe > .aBBjbd { animation: 0.3s ease-out 0s 1 normal forwards running quantumWizBoxInkSpread; background-image: radial-gradient(circle farthest-side, rgb(189, 189, 189), rgb(189, 189, 189) 80%, rgba(189, 189, 189, 0) 100%); background-size: cover; opacity: 1; top: 0px; left: 0px; }

.J0XlZe { color: inherit; line-height: 40px; padding: 0px 6px 0px 1em; }

.a9caSc { color: inherit; direction: ltr; padding: 0px 6px 0px 1em; }

.kCtYwe { border-top: 1px solid rgba(0, 0, 0, 0.12); margin: 7px 0px; }

.B2l7lc { border-left: 1px solid rgba(0, 0, 0, 0.12); display: inline-block; height: 48px; }

@media screen and (max-width: 840px) {
  .JAPqpe { padding: 8px 0px; }
  .z80M1 { padding: 0px 16px; }
  .JPdR6b.e5Emjc .z80M1 { padding-left: 48px; }
  .PCdOIb { left: 12px; }
}

.oxMpi { padding: 0px 16px 18px; }

.hB0k6, .ZtDwgb { margin-right: 8px; }

.hB0k6, .QX73N, .ZtDwgb { padding: 0px 16px; }

.hB0k6, .QX73N { border-radius: var(--dt-corner-button,.25rem); }

.AOYJ6c { height: 48px; width: 100%; }

.AOYJ6c, .AOYJ6c .VfPpkd-Jh9lGc { border-radius: 100px; }

.oxMpi .AOYJ6c .MaxOIc { font-size: 24px; height: 24px; width: 24px; }

.SSMtpf { font: var(--dt-label-small-font,500 .6875rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-small-spacing,.0727272727em); text-transform: var(--dt-label-small-transform,uppercase); color: var(--dt-on-surface,rgb(60,64,67)); padding-bottom: 16px; }

.TUd9Hf { display: flex; -webkit-box-flex: 1; flex: 1 1 auto; margin-bottom: 14px; }

.aKBAzc { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.ah4wbe { -webkit-box-flex: 1; flex: 1 1 auto; word-break: break-word; }

.Rz1NYe { display: flex; padding-bottom: 12px; }

.aCNyvf { padding-right: 14px; }

.j5TJQ { font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,.0178571429em); color: var(--dt-on-surface,rgb(60,64,67)); }

.jtn0Vb { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); color: var(--dt-on-surface,rgb(60,64,67)); user-select: text; white-space: pre-line; }

.AYfYVc, .s2aAtd { padding-top: 4px; }

.m99ddd, .xt4Y1d { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); color: var(--dt-on-surface,rgb(60,64,67)); }

.Rz1NYe .m99ddd { font-weight: 400; }

.J3TqDb, .nhkJid, .QYAGmd { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); color: var(--dt-on-surface,rgb(60,64,67)); padding-bottom: 4px; }

.hiEOsf, .PHm6qf { display: flex; -webkit-box-flex: 1; flex-grow: 1; font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); }

.hiEOsf { color: var(--dt-on-surface,rgb(60,64,67)); }

.PHm6qf { color: var(--dt-on-surface-variant,rgb(95,99,104)); text-decoration: line-through; }

.Dw6xSd { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); color: var(--dt-on-surface,rgb(60,64,67)); }

.Z58F5b { color: var(--dt-tertiary,rgb(24,128,56)); }

.YuNKGb { color: var(--dt-error,rgb(217,48,37)); }

.BQynZe { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.cKL5M { height: 35px; width: 35px; }

.lPQaNe .If2P7d { border: none; display: flex; margin-bottom: 16px; -webkit-box-orient: vertical; -webkit-box-direction: reverse; flex-direction: column-reverse; }

.lPQaNe .GMQ90d { border: none; padding: 0px; margin: 0px; }

.BOcHJe { -webkit-box-align: center; align-items: center; display: flex; width: 100%; }

.vehxkc { -webkit-box-align: stretch; align-items: stretch; border: 1px solid rgba(0, 0, 0, 0.08); border-radius: 4px; display: flex; -webkit-box-pack: justify; justify-content: space-between; margin: 14px; padding: 3px 6px 3px 10px; }

.BEmwVc { border-top: 1px solid rgba(0, 0, 0, 0.08); }

.j1UHoe { display: none; padding: 2px; }

.j1UHoe .FMvKQd { margin-top: 0px; }

.BEmwVc.rmm4Cf .O0NXze { display: none; }

.BEmwVc.rmm4Cf .j1UHoe { display: block; }

.O0NXze { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: end; justify-content: flex-end; margin: 0px -0.5rem 0px 0.25rem; padding: 0px; }

.O0NXze .VfPpkd-kBDsod { display: flex; }

.vFuuxf { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; margin-right: -2px; -webkit-box-pack: end; justify-content: flex-end; }

.vFuuxf .O0NXze .HXRT5b { height: 24px; width: 24px; }

.edhGSc { user-select: none; -webkit-tap-highlight-color: transparent; display: inline-block; outline: none; padding-bottom: 8px; }

.RpC4Ne { min-height: 1.5em; position: relative; vertical-align: top; }

.Pc9Gce { display: flex; position: relative; padding-top: 14px; }

.KHxj8b { -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; background-color: transparent; border: none; display: block; font: 400 16px / 24px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 24px; min-height: 24px; margin: 0px; outline: none; padding: 0px; resize: none; white-space: pre-wrap; overflow-wrap: break-word; z-index: 0; overflow: hidden visible; }

.KHxj8b.VhWN2c { text-align: center; }

.edhGSc.dm7YTc .KHxj8b { color: rgba(255, 255, 255, 0.87); }

.edhGSc.u3bW4e.dm7YTc .KHxj8b { color: rgb(255, 255, 255); }

.z0oSpf { background-color: rgba(0, 0, 0, 0.12); height: 1px; left: 0px; margin: 0px; padding: 0px; position: absolute; width: 100%; }

.edhGSc.dm7YTc > .RpC4Ne > .z0oSpf { background-color: rgba(255, 255, 255, 0.12); }

.Bfurwb { transform: scaleX(0); background-color: rgb(66, 133, 244); height: 2px; left: 0px; margin: 0px; padding: 0px; position: absolute; width: 100%; }

.edhGSc.k0tWj > .RpC4Ne > .z0oSpf, .edhGSc.k0tWj > .RpC4Ne > .Bfurwb { background-color: rgb(213, 0, 0); height: 2px; }

.edhGSc.k0tWj.dm7YTc > .RpC4Ne > .z0oSpf, .edhGSc.k0tWj.dm7YTc > .RpC4Ne > .Bfurwb { background-color: rgb(255, 110, 110); }

.edhGSc.RDPZE .KHxj8b { color: rgba(0, 0, 0, 0.38); }

.edhGSc.RDPZE > .RpC4Ne > .z0oSpf { background: none; border-bottom: 1px dotted rgba(0, 0, 0, 0.38); }

.Bfurwb.Y2Zypf { animation: 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running quantumWizPaperInputRemoveUnderline; }

.edhGSc.u3bW4e > .RpC4Ne > .Bfurwb { animation: 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running quantumWizPaperInputAddUnderline; transform: scaleX(1); }

.edhGSc.FPYHkb > .RpC4Ne { padding-top: 24px; }

.fqp6hd { transform-origin: left top; transform: translate(0px, -22px); transition: color 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s, top, transform, -webkit-transform; color: rgba(0, 0, 0, 0.38); font: 400 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; pointer-events: none; position: absolute; top: 100%; width: 100%; }

.edhGSc.u3bW4e > .RpC4Ne > .fqp6hd, .edhGSc.CDELXb > .RpC4Ne > .fqp6hd, .edhGSc.LydCob .fqp6hd { transform: scale(0.75); top: 16px; }

.edhGSc.dm7YTc > .RpC4Ne > .fqp6hd { color: rgba(255, 255, 255, 0.38); }

.edhGSc.u3bW4e > .RpC4Ne > .fqp6hd, .edhGSc.u3bW4e.dm7YTc > .RpC4Ne > .fqp6hd { color: rgb(66, 133, 244); }

.F1pOBe { color: rgba(0, 0, 0, 0.38); font: 400 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; max-width: 100%; overflow: hidden; pointer-events: none; position: absolute; bottom: 3px; text-overflow: ellipsis; white-space: nowrap; }

.edhGSc.dm7YTc .F1pOBe { color: rgba(255, 255, 255, 0.38); }

.edhGSc.CDELXb > .RpC4Ne > .F1pOBe { display: none; }

.S1BUyf { -webkit-tap-highlight-color: transparent; font: 400 12px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 16px; margin-left: auto; padding-left: 16px; padding-top: 8px; pointer-events: none; text-align: right; color: rgba(0, 0, 0, 0.38); white-space: nowrap; }

.edhGSc.dm7YTc > .S1BUyf { color: rgba(255, 255, 255, 0.38); }

.edhGSc.wrxyb { padding-bottom: 4px; }

.v6odTb, .YElZX:not(:empty) { -webkit-tap-highlight-color: transparent; -webkit-box-flex: 1; flex: 1 1 auto; font: 400 12px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; min-height: 16px; padding-top: 8px; }

.edhGSc.wrxyb .jE8NUc { display: flex; }

.YElZX { pointer-events: none; }

.v6odTb { color: rgb(213, 0, 0); }

.edhGSc.dm7YTc .v6odTb { color: rgb(255, 110, 110); }

.YElZX { opacity: 0.3; }

.edhGSc.k0tWj .YElZX, .edhGSc:not(.k0tWj) .YElZX:not(:empty) + .v6odTb { display: none; }

@-webkit-keyframes quantumWizPaperInputRemoveUnderline { 
  0% { transform: scaleX(1); opacity: 1; }
  100% { transform: scaleX(1); opacity: 0; }
}

@keyframes quantumWizPaperInputRemoveUnderline { 
  0% { transform: scaleX(1); opacity: 1; }
  100% { transform: scaleX(1); opacity: 0; }
}

@-webkit-keyframes quantumWizPaperInputAddUnderline { 
  0% { transform: scaleX(0); }
  100% { transform: scaleX(1); }
}

@keyframes quantumWizPaperInputAddUnderline { 
  0% { transform: scaleX(0); }
  100% { transform: scaleX(1); }
}

.ZAJxef, .eYTr6c { height: 32px; position: relative; width: 32px; }

.LZ2FEb { animation: 0.27s linear 0s 1 normal backwards running animateApprovalPersonIconIn; border-radius: 50%; height: 32px; opacity: 1; width: 32px; }

@-webkit-keyframes animateApprovalPersonIconIn { 
  0% { opacity: 0; }
}

@keyframes animateApprovalPersonIconIn { 
  0% { opacity: 0; }
}

.oJg3bc, .IXkYsf, .OGF2Yc { height: 20px; position: relative; width: 20px; }

.OGF2Yc { border-radius: 50%; }

.ZAJxef, .oJg3bc { display: inline-flex; }

.eYTr6c { border-radius: 16px; background-color: var(--dt-surface-variant,rgb(241,243,244)); }

.IXkYsf { border-radius: 10px; }

.Kjmrtb { left: 24px; position: absolute; top: 20px; }

.lxuawb { background-color: var(--dt-surface2,#fff); border-radius: 50%; height: 18px; position: absolute; width: 18px; }

.zX4kg { border-radius: var(--dt-corner-landmark,0); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow-y: auto; }

.cKrIre { height: 100vh; max-width: 320px; }

.FSIBbb { -webkit-box-align: center; align-items: center; display: flex; height: 64px; margin: 1px; -webkit-box-pack: justify; justify-content: space-between; }

.zjwBT { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.MX9Vje { display: flex; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; }

.oW88wd { position: relative; }

.Ag6gR { font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,.00625em); color: var(--dt-on-surface,rgb(60,64,67)); display: flex; -webkit-box-flex: 1; flex: 1 1 auto; }

.CS5vN { color: var(--dt-primary,rgb(26,115,232)); margin-right: 20px; vertical-align: middle; }

.hATPff { display: flex; -webkit-box-flex: 1; flex: 1 1 auto; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; height: 93%; overflow-y: auto; }

.BtuWMb .hATPff { display: flex; overflow-y: auto; }

.siStgd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 auto; }

.xEacub .QIrpef, .DPnoGc .QIrpef { color: var(--dt-on-surface-variant,rgb(95,99,104)); height: 1.25rem; width: 1.25rem; }

.B8vHne { fill: var(--dt-on-surface-variant,rgb(95,99,104)); }

.BtuWMb .ncWkde { fill: var(--dt-primary-container-icon,rgb(25,103,210)); }

.BtuWMb .wJZ8Wb .gGYsWb { color: var(--dt-primary-action,rgb(25,103,210)); }

.BtuWMb .wJZ8Wb .gGYsWb, .BtuWMb .wJZ8Wb .gGYsWb::before, .BtuWMb .wJZ8Wb .gGYsWb::after { background-color: var(--dt-primary-container,rgb(232,240,254)); }

.DPnoGc { position: absolute; top: 10px; }

.wP8nMd { border-top: solid 1px var(--dt-outline-variant,rgb(218,220,224)); }

.olFVe { padding-left: 8px; }

.olFVe .M26Hse { height: 35px; padding: 0px 8px; }

.A4y5Eb { padding: 0px 15px 18px; }

.H7Syve { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: justify; justify-content: space-between; }

.B3P4Pe { color: var(--dt-on-surface,rgb(60,64,67)); font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-stretch: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; text-transform: var(--dt-label-small-transform,uppercase); font-size: 11px; font-weight: 500; letter-spacing: 0.4px; padding-bottom: 8px; }

.nh7RAf { height: 375px; }

.siStgd .nh7RAf .If2P7d { display: none; }

.UmQeIf { -webkit-box-align: center; align-items: center; background-color: var(--dt-scrim,rgba(32,33,36,.6)); display: flex; position: absolute; height: 100%; width: 100%; z-index: 1; }

.ysbVIc { margin-top: 0px; }

.sBvv3 { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; }

.J0Td4b { -webkit-box-align: center; align-items: center; display: flex; }

.RpcR8e { border-top: 1px solid var(--dt-outline-variant,rgb(218,220,224)); margin: 0px 15px 10px; }

.A30Pgc { border-radius: 8px; left: 50%; top: 50%; transform: translateX(-50%) translateY(-50%); }

.L0UvRd { width: 100%; }

.i6N7Re .qFjdb.JV458b { color: var(--dt-error,rgb(217,48,37)); fill: currentcolor; }

.i6N7Re .qFjdb.do04jc { color: var(--dt-tertiary,rgb(24,128,56)); fill: currentcolor; }

.i6N7Re .qFjdb.S42Ve { color: var(--dt-primary-action,rgb(25,103,210)); fill: currentcolor; }

.i6N7Re { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; padding: 16px 16px 14px 20px; }

.FvWGJd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex-grow: 1; }

.WGUH5e { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); padding-top: 4px; }

.pHw1O { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.ZhJ4ge .FvWGJd { padding-left: 200px; }

.x1pG1e { font: var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-large-spacing,0); -webkit-box-flex: 1; flex-grow: 1; }

.tnFpPb { height: 48px; margin-bottom: -4px; padding-top: 4px; width: auto; }

.gUU7vb { color: var(--dt-on-surface-variant,rgb(95,99,104)); margin-right: -12px; }

.P6msMd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 auto; padding: 0px 15px; }

.P6msMd.LsH4n { -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-pack: justify; justify-content: space-between; overflow-y: auto; }

.BCOcpf { display: flex; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: justify; justify-content: space-between; }

.LsH4n .BCOcpf { padding-right: 30px; width: 170px; }

.ne9O6d { -webkit-box-flex: 0; flex: 0 0 auto; padding-bottom: 15px; }

.tWS7Jd { min-height: 44px; }

.xAev4e { -webkit-box-flex: 1; flex: 1 1 auto; min-height: 200px; }

.oBIJVb { -webkit-box-align: center; align-items: center; display: flex; height: 48px; -webkit-box-pack: justify; justify-content: space-between; }

.V24RSd .oBIJVb { -webkit-box-align: baseline; align-items: baseline; height: 32px; }

.SKM7kf { color: var(--dt-on-surface,rgb(60,64,67)); margin-right: -12px; }

.vRUySd { font: var(--dt-label-medium-font,500 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-medium-spacing,.0208333333em); color: var(--dt-primary-container-link,rgb(25,103,210)); display: inline-block; margin: 12px 0px 16px; }

.Zsj9Fd { color: var(--dt-on-surface,rgb(60,64,67)); font: var(--dt-label-small-font,500 .6875rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-small-spacing,.0727272727em); text-transform: var(--dt-label-small-transform,uppercase); }

.tIgSeb { display: flex; justify-self: flex-start; min-height: 50px; }

.V24RSd .srcFDf { padding-bottom: 0px; }

.srcFDf { padding-bottom: 16px; }

.yLLlPc { padding-right: 16px; }

.emszSc { color: var(--dt-on-surface,rgb(60,64,67)); max-width: 150px; overflow: hidden; text-overflow: ellipsis; font: var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-label-large-spacing,.0178571429em); }

.boO95 { color: var(--dt-on-surface-variant,rgb(95,99,104)); font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); }

.AjmcOb { padding-left: 8px; }

.tJhwNb { color: var(--dt-on-surface-variant,rgb(95,99,104)); margin-left: auto; margin-right: -8px; }

.PYrZc { width: inherit; }

.UqvRcc { box-sizing: border-box; display: inline-block; position: relative; max-height: 100%; max-width: 100%; width: inherit; }

.VrQwO { display: none; }

.sbsxqb { pointer-events: none; transition: opacity 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0.15s; inset: 0px; position: fixed; opacity: 0; z-index: 5000; background-color: rgba(0, 0, 0, 0.5); }

.sbsxqb.iWO5td { pointer-events: all; transition: opacity 0.05s cubic-bezier(0.4, 0, 0.2, 1) 0s; opacity: 1; }

@-webkit-keyframes primary-indeterminate-translate { 
  0% { transform: translateX(-145.167%); }
  20% { animation-timing-function: cubic-bezier(0.5, 0, 0.701732, 0.495819); transform: translateX(-145.167%); }
  59.15% { animation-timing-function: cubic-bezier(0.302435, 0.381352, 0.55, 0.956352); transform: translateX(-61.4952%); }
  100% { transform: translateX(55.4444%); }
}

@keyframes primary-indeterminate-translate { 
  0% { transform: translateX(-145.167%); }
  20% { animation-timing-function: cubic-bezier(0.5, 0, 0.701732, 0.495819); transform: translateX(-145.167%); }
  59.15% { animation-timing-function: cubic-bezier(0.302435, 0.381352, 0.55, 0.956352); transform: translateX(-61.4952%); }
  100% { transform: translateX(55.4444%); }
}

@-webkit-keyframes primary-indeterminate-translate-reverse { 
  0% { transform: translateX(145.167%); }
  20% { animation-timing-function: cubic-bezier(0.5, 0, 0.701732, 0.495819); transform: translateX(145.167%); }
  59.15% { animation-timing-function: cubic-bezier(0.302435, 0.381352, 0.55, 0.956352); transform: translateX(61.4952%); }
  100% { transform: translateX(-55.4444%); }
}

@keyframes primary-indeterminate-translate-reverse { 
  0% { transform: translateX(145.167%); }
  20% { animation-timing-function: cubic-bezier(0.5, 0, 0.701732, 0.495819); transform: translateX(145.167%); }
  59.15% { animation-timing-function: cubic-bezier(0.302435, 0.381352, 0.55, 0.956352); transform: translateX(61.4952%); }
  100% { transform: translateX(-55.4444%); }
}

@-webkit-keyframes primary-indeterminate-scale { 
  0% { transform: scaleX(0.08); }
  36.65% { animation-timing-function: cubic-bezier(0.334731, 0.12482, 0.785844, 1); transform: scaleX(0.08); }
  69.15% { animation-timing-function: cubic-bezier(0.06, 0.11, 0.6, 1); transform: scaleX(0.661479); }
  100% { transform: scaleX(0.08); }
}

@keyframes primary-indeterminate-scale { 
  0% { transform: scaleX(0.08); }
  36.65% { animation-timing-function: cubic-bezier(0.334731, 0.12482, 0.785844, 1); transform: scaleX(0.08); }
  69.15% { animation-timing-function: cubic-bezier(0.06, 0.11, 0.6, 1); transform: scaleX(0.661479); }
  100% { transform: scaleX(0.08); }
}

@-webkit-keyframes auxiliary-indeterminate-translate { 
  0% { animation-timing-function: cubic-bezier(0.15, 0, 0.515058, 0.409685); transform: translateX(-54.8889%); }
  25% { animation-timing-function: cubic-bezier(0.31033, 0.284058, 0.8, 0.733712); transform: translateX(-17.237%); }
  48.35% { animation-timing-function: cubic-bezier(0.4, 0.627035, 0.6, 0.902026); transform: translateX(29.4973%); }
  100% { transform: translateX(105.389%); }
}

@keyframes auxiliary-indeterminate-translate { 
  0% { animation-timing-function: cubic-bezier(0.15, 0, 0.515058, 0.409685); transform: translateX(-54.8889%); }
  25% { animation-timing-function: cubic-bezier(0.31033, 0.284058, 0.8, 0.733712); transform: translateX(-17.237%); }
  48.35% { animation-timing-function: cubic-bezier(0.4, 0.627035, 0.6, 0.902026); transform: translateX(29.4973%); }
  100% { transform: translateX(105.389%); }
}

@-webkit-keyframes auxiliary-indeterminate-translate-reverse { 
  0% { animation-timing-function: cubic-bezier(0.15, 0, 0.515058, 0.409685); transform: translateX(54.8889%); }
  25% { animation-timing-function: cubic-bezier(0.31033, 0.284058, 0.8, 0.733712); transform: translateX(17.237%); }
  48.35% { animation-timing-function: cubic-bezier(0.4, 0.627035, 0.6, 0.902026); transform: translateX(-29.4973%); }
  100% { transform: translateX(-105.389%); }
}

@keyframes auxiliary-indeterminate-translate-reverse { 
  0% { animation-timing-function: cubic-bezier(0.15, 0, 0.515058, 0.409685); transform: translateX(54.8889%); }
  25% { animation-timing-function: cubic-bezier(0.31033, 0.284058, 0.8, 0.733712); transform: translateX(17.237%); }
  48.35% { animation-timing-function: cubic-bezier(0.4, 0.627035, 0.6, 0.902026); transform: translateX(-29.4973%); }
  100% { transform: translateX(-105.389%); }
}

@-webkit-keyframes auxiliary-indeterminate-scale { 
  0% { animation-timing-function: cubic-bezier(0.205028, 0.057051, 0.57661, 0.453971); transform: scaleX(0.08); }
  19.15% { animation-timing-function: cubic-bezier(0.152313, 0.196432, 0.648374, 1.00432); transform: scaleX(0.457104); }
  44.15% { animation-timing-function: cubic-bezier(0.257759, 0.003163, 0.211762, 1.38179); transform: scaleX(0.72796); }
  100% { transform: scaleX(0.08); }
}

@keyframes auxiliary-indeterminate-scale { 
  0% { animation-timing-function: cubic-bezier(0.205028, 0.057051, 0.57661, 0.453971); transform: scaleX(0.08); }
  19.15% { animation-timing-function: cubic-bezier(0.152313, 0.196432, 0.648374, 1.00432); transform: scaleX(0.457104); }
  44.15% { animation-timing-function: cubic-bezier(0.257759, 0.003163, 0.211762, 1.38179); transform: scaleX(0.72796); }
  100% { transform: scaleX(0.08); }
}

@-webkit-keyframes buffering { 
  100% { transform: translateX(-10px); }
}

@keyframes buffering { 
  100% { transform: translateX(-10px); }
}

@-webkit-keyframes buffering-reverse { 
  100% { transform: translateX(10px); }
}

@keyframes buffering-reverse { 
  100% { transform: translateX(10px); }
}

@-webkit-keyframes indeterminate-translate-ie { 
  0% { transform: translateX(-100%); }
  100% { transform: translateX(100%); }
}

@keyframes indeterminate-translate-ie { 
  0% { transform: translateX(-100%); }
  100% { transform: translateX(100%); }
}

@-webkit-keyframes indeterminate-translate-reverse-ie { 
  0% { transform: translateX(100%); }
  100% { transform: translateX(-100%); }
}

@keyframes indeterminate-translate-reverse-ie { 
  0% { transform: translateX(100%); }
  100% { transform: translateX(-100%); }
}

.sZwd7c { height: 4px; overflow: hidden; position: relative; transform: translateZ(0px); transition: opacity 250ms linear 0s; width: 100%; }

.w2zcLc { position: absolute; }

.xcNBHc, .MyvhI, .l3q5xe { height: 100%; position: absolute; width: 100%; }

.w2zcLc { transform-origin: left top; transition: transform 250ms ease 0s, -webkit-transform 250ms ease 0s; }

.MyvhI { transform-origin: left top; transition: transform 250ms ease 0s, -webkit-transform 250ms ease 0s; animation: 0s ease 0s 1 normal none running none; }

.l3q5xe { animation: 0s ease 0s 1 normal none running none; }

.w2zcLc { background-color: rgb(230, 230, 230); height: 100%; transform-origin: left top; transition: transform 250ms ease 0s, -webkit-transform 250ms ease 0s; width: 100%; }

.TKVRUb { transform: scaleX(0); }

.sUoeld { visibility: hidden; }

.l3q5xe { background-color: rgb(0, 0, 0); display: inline-block; }

.xcNBHc { background-size: 10px 4px; background-repeat: repeat-x; background-image: url("data:image/svg+xml;charset=UTF-8,%3Csvg%20version%3D%271.1%27%20xmlns%3D%27http%3A%2F%2Fwww.w3.org%2F2000%2Fsvg%27%20xmlns%3Axlink%3D%27http%3A%2F%2Fwww.w3.org%2F1999%2Fxlink%27%20x%3D%270px%27%20y%3D%270px%27%20enable-background%3D%27new%200%200%205%202%27%20xml%3Aspace%3D%27preserve%27%20viewBox%3D%270%200%205%202%27%20preserveAspectRatio%3D%27none%20slice%27%3E%3Ccircle%20cx%3D%271%27%20cy%3D%271%27%20r%3D%271%27%20fill%3D%27%23e6e6e6%27%2F%3E%3C%2Fsvg%3E"); visibility: hidden; }

.sZwd7c.B6Vhqe .MyvhI { transition: none 0s ease 0s; }

.sZwd7c.B6Vhqe .TKVRUb { animation: 2s linear 0s infinite normal none running primary-indeterminate-translate; }

.sZwd7c.B6Vhqe .TKVRUb > .l3q5xe { animation: 2s linear 0s infinite normal none running primary-indeterminate-scale; }

.sZwd7c.B6Vhqe .sUoeld { animation: 2s linear 0s infinite normal none running auxiliary-indeterminate-translate; visibility: visible; }

.sZwd7c.B6Vhqe .sUoeld > .l3q5xe { animation: 2s linear 0s infinite normal none running auxiliary-indeterminate-scale; }

.sZwd7c.B6Vhqe.ieri7c .l3q5xe { transform: scaleX(0.45); }

.sZwd7c.B6Vhqe.ieri7c .sUoeld { animation: 0s ease 0s 1 normal none running none; visibility: hidden; }

.sZwd7c.B6Vhqe.ieri7c .TKVRUb { animation: 2s ease-out 0s infinite normal none running indeterminate-translate-ie; }

.sZwd7c.B6Vhqe.ieri7c .TKVRUb > .l3q5xe, .sZwd7c.B6Vhqe.ieri7c .sUoeld > .l3q5xe { animation: 0s ease 0s 1 normal none running none; }

.sZwd7c.juhVM .w2zcLc, .sZwd7c.juhVM .MyvhI { right: 0px; transform-origin: right center; }

.sZwd7c.juhVM .TKVRUb { animation-name: primary-indeterminate-translate-reverse; }

.sZwd7c.juhVM .sUoeld { animation-name: auxiliary-indeterminate-translate-reverse; }

.sZwd7c.juhVM.ieri7c .TKVRUb { animation-name: indeterminate-translate-reverse-ie; }

.sZwd7c.qdulke { opacity: 0; }

.sZwd7c.jK7moc .sUoeld, .sZwd7c.jK7moc .TKVRUb, .sZwd7c.jK7moc .sUoeld > .l3q5xe, .sZwd7c.jK7moc .TKVRUb > .l3q5xe { animation-play-state: paused; }

.sZwd7c.D6TUi .xcNBHc { animation: 250ms linear 0s infinite normal none running buffering; visibility: visible; }

.sZwd7c.D6TUi.juhVM .xcNBHc { animation: 250ms linear 0s infinite normal none running buffering-reverse; }

.RM9ulf { visibility: hidden; position: fixed; z-index: 5000; color: rgb(255, 255, 255); pointer-events: none; }

.RM9ulf.catR2e { max-width: 90%; max-height: 90%; }

.R8qYlc { border-radius: 2px; background-color: rgba(97, 97, 97, 0.9); position: absolute; left: 0px; width: 100%; height: 100%; opacity: 0; transform: scale(0, 0.5); transform-origin: inherit; }

.AZnilc { display: block; position: relative; font-size: 10px; font-weight: 500; padding: 5px 8px 6px; opacity: 0; }

.RM9ulf.qs41qe .R8qYlc { opacity: 1; transform: scale(1, 1); }

.RM9ulf.catR2e .AZnilc { overflow-wrap: break-word; }

.RM9ulf.qs41qe .AZnilc { opacity: 1; }

.RM9ulf.AXm5jc .AZnilc { font-size: 14px; padding: 8px 16px; }

.RM9ulf.u5lFJe { transition-property: transform, -webkit-transform; transition-duration: 200ms; transition-timing-function: cubic-bezier(0.24, 1, 0.32, 1); }

.RM9ulf.u5lFJe .R8qYlc { transition-property: opacity, transform, -webkit-transform; transition-duration: 50ms, 200ms; transition-timing-function: linear, cubic-bezier(0.24, 1, 0.32, 1); }

.RM9ulf.u5lFJe .AZnilc { transition: opacity 150ms cubic-bezier(0, 0, 0.6, 1) 50ms; }

.RM9ulf.xCxor { transition: opacity 70ms linear 0ms; }

.O0WRkf { user-select: none; transition: background 0.2s ease 0.1s; border: 0px; border-radius: 3px; cursor: pointer; display: inline-block; font-size: 14px; font-weight: 500; min-width: 4em; outline: none; overflow: hidden; position: relative; text-align: center; text-transform: uppercase; -webkit-tap-highlight-color: transparent; z-index: 0; }

.A9jyad { font-size: 13px; line-height: 16px; }

.zZhnYe { transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; background: rgb(223, 223, 223); box-shadow: rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 3px 1px -2px, rgba(0, 0, 0, 0.2) 0px 1px 5px 0px; }

.zZhnYe.qs41qe { transition: background 0.8s ease 0s; box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; }

.e3Duub, .e3Duub a, .e3Duub a:hover, .e3Duub a:link, .e3Duub a:visited { background: rgb(66, 133, 244); color: rgb(255, 255, 255); }

.HQ8yf, .HQ8yf a { color: rgb(66, 133, 244); }

.UxubU, .UxubU a { color: rgb(255, 255, 255); }

.ZFr60d { position: absolute; inset: 0px; background-color: transparent; }

.O0WRkf.u3bW4e .ZFr60d { background-color: rgba(0, 0, 0, 0.12); }

.UxubU.u3bW4e .ZFr60d { background-color: rgba(255, 255, 255, 0.3); }

.e3Duub.u3bW4e .ZFr60d { background-color: rgba(0, 0, 0, 0.12); }

.HQ8yf.u3bW4e .ZFr60d { background-color: rgba(66, 133, 244, 0.15); }

.Vwe4Vb { transform: translate(-50%, -50%) scale(0); transition: opacity 0.2s ease 0s, visibility 0s ease 0.2s, -webkit-transform 0s ease 0.2s; background-size: cover; left: 0px; opacity: 0; pointer-events: none; position: absolute; top: 0px; visibility: hidden; }

.O0WRkf.qs41qe .Vwe4Vb { transform: translate(-50%, -50%) scale(2.2); opacity: 1; visibility: visible; }

.O0WRkf.qs41qe.M9Bg4d .Vwe4Vb { transition: transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s, opacity 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, -webkit-transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s; }

.O0WRkf.j7nIZb .Vwe4Vb { transform: translate(-50%, -50%) scale(2.2); visibility: visible; }

.oG5Srb .Vwe4Vb, .zZhnYe .Vwe4Vb { background-image: radial-gradient(circle farthest-side, rgba(0, 0, 0, 0.12), rgba(0, 0, 0, 0.12) 80%, rgba(0, 0, 0, 0) 100%); }

.HQ8yf .Vwe4Vb { background-image: radial-gradient(circle farthest-side, rgba(66, 133, 244, 0.25), rgba(66, 133, 244, 0.25) 80%, rgba(66, 133, 244, 0) 100%); }

.e3Duub .Vwe4Vb { background-image: radial-gradient(circle farthest-side, rgb(51, 103, 214), rgb(51, 103, 214) 80%, rgba(51, 103, 214, 0) 100%); }

.UxubU .Vwe4Vb { background-image: radial-gradient(circle farthest-side, rgba(255, 255, 255, 0.3), rgba(255, 255, 255, 0.3) 80%, rgba(255, 255, 255, 0) 100%); }

.O0WRkf.RDPZE { box-shadow: none; color: rgba(68, 68, 68, 0.5); cursor: default; fill: rgba(68, 68, 68, 0.5); }

.zZhnYe.RDPZE { background: rgba(153, 153, 153, 0.1); }

.UxubU.RDPZE { color: rgba(255, 255, 255, 0.5); fill: rgba(255, 255, 255, 0.5); }

.UxubU.zZhnYe.RDPZE { background: rgba(204, 204, 204, 0.1); }

.CwaK9 { position: relative; }

.RveJvd { display: inline-block; margin: 0.5em; }

.XHsn7e { background-color: rgb(0, 0, 0); border: none; border-radius: 50%; box-sizing: content-box; box-shadow: rgba(0, 0, 0, 0.14) 0px 6px 10px 0px, rgba(0, 0, 0, 0.12) 0px 1px 18px 0px, rgba(0, 0, 0, 0.2) 0px 3px 5px -1px; cursor: pointer; display: inline-block; fill: rgb(255, 255, 255); height: 56px; outline: none; overflow: hidden; position: relative; text-align: center; width: 56px; z-index: 4000; }

.HaXdpb { background: rgba(255, 255, 255, 0.2); inset: 0px; display: none; position: absolute; }

.XHsn7e:hover { box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; }

.XHsn7e:hover .HaXdpb { display: block; }

.XHsn7e.qs41qe { box-shadow: rgba(0, 0, 0, 0.14) 0px 12px 17px 2px, rgba(0, 0, 0, 0.12) 0px 5px 22px 4px, rgba(0, 0, 0, 0.2) 0px 7px 8px -4px; }

.XHsn7e.qs41qe .HaXdpb { display: block; }

.XHsn7e.RDPZE { background: rgba(153, 153, 153, 0.1); box-shadow: none; color: rgba(68, 68, 68, 0.5); cursor: default; fill: rgba(68, 68, 68, 0.5); }

.XHsn7e.RDPZE:hover { opacity: 1; }

.XHsn7e.RDPZE .HaXdpb { display: none; }

.XHsn7e:focus { box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; }

.XHsn7e:focus .HaXdpb { display: block; }

.Ip8zfc { display: inline-block; height: 24px; position: absolute; top: 16px; left: 16px; width: 24px; transform: rotate(0deg); transition: all 0.3s ease-in-out 0s; }

.Ip8zfc.eLNT1d { opacity: 0; visibility: hidden; transform: rotate(225deg); transition: all 0.3s ease-in-out 0s; }

.Ip8zfc.ReqAjb { transform: rotate(135deg); transition: all 0.3s ease-in-out 0s; }

.dURtfb { height: 40px; width: 40px; }

.dURtfb .Ip8zfc { top: 8px; left: 8px; }

.HRp7vf { transform: translate(-50%, -50%) scale(0); transition: opacity 0.2s ease 0s, visibility 0s ease 0.2s, -webkit-transform 0s ease 0.2s; background-image: radial-gradient(circle farthest-side, rgba(204, 204, 204, 0.25), rgba(204, 204, 204, 0.25) 80%, rgba(204, 204, 204, 0) 100%); background-size: cover; left: 0px; opacity: 0; pointer-events: none; position: absolute; top: 0px; visibility: hidden; }

.XHsn7e.qs41qe > .HRp7vf { transform: translate(-50%, -50%) scale(2.2); opacity: 1; visibility: visible; }

.XHsn7e.qs41qe.M9Bg4d > .HRp7vf { transition: transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s, opacity 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, -webkit-transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s; }

.XHsn7e.j7nIZb > .HRp7vf { transform: translate(-50%, -50%) scale(2.2); visibility: visible; }

.cTPETe { display: flex; }

.u1Djpb { display: flex; height: 22px; border-radius: 11px; margin: 0px 6px 0px 0px; padding-left: 12px; white-space: nowrap; color: rgba(0, 0, 0, 0.87); background-color: rgb(224, 224, 224); font-size: 14px; }

.fb31zf { margin: auto; }

.GorKAf { display: inline-block; position: relative; margin: 3px; width: 16px; height: 16px; background-color: rgba(0, 0, 0, 0.38); border-radius: 50%; }

.GorKAf::before, .GorKAf::after { content: ""; position: absolute; width: 10px; height: 2px; top: 7px; background-color: rgb(224, 224, 224); }

.GorKAf::before { transform: rotate(45deg); left: 3px; }

.GorKAf::after { transform: rotate(-45deg); right: 3px; }

.u1Djpb:hover { color: white; }

.u1Djpb:hover, .u1Djpb:hover .GorKAf::before, .u1Djpb:hover .GorKAf::after { background-color: rgb(97, 97, 97); }

.u1Djpb:hover .GorKAf { background-color: white; }

.rFrNMe { user-select: none; -webkit-tap-highlight-color: transparent; display: inline-block; outline: none; padding-bottom: 8px; width: 200px; }

.aCsJod { height: 40px; position: relative; vertical-align: top; }

.aXBtI { display: flex; position: relative; top: 14px; }

.Xb9hP { display: flex; -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; min-width: 0%; position: relative; }

.A37UZe { box-sizing: border-box; height: 24px; line-height: 24px; position: relative; }

.qgcB3c:not(:empty) { padding-right: 12px; }

.sxyYjd:not(:empty) { padding-left: 12px; }

.whsOnd { -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; background-color: transparent; border: none; display: block; font: 400 16px / 24px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 24px; margin: 0px; min-width: 0%; outline: none; padding: 0px; z-index: 0; }

.rFrNMe.dm7YTc .whsOnd { color: rgb(255, 255, 255); }

.i9lrp { background-color: rgba(0, 0, 0, 0.12); bottom: -2px; height: 1px; left: 0px; margin: 0px; padding: 0px; position: absolute; width: 100%; }

.i9lrp::before { content: ""; position: absolute; inset: 0px 0px -2px; border-bottom: 1px solid rgba(0, 0, 0, 0); pointer-events: none; }

.rFrNMe.dm7YTc .i9lrp { background-color: rgba(255, 255, 255, 0.7); }

.OabDMe { transform: scaleX(0); background-color: rgb(66, 133, 244); bottom: -2px; height: 2px; left: 0px; margin: 0px; padding: 0px; position: absolute; width: 100%; }

.rFrNMe.dm7YTc .OabDMe { background-color: rgb(161, 194, 250); }

.rFrNMe.k0tWj .i9lrp, .rFrNMe.k0tWj .OabDMe { background-color: rgb(213, 0, 0); height: 2px; }

.rFrNMe.k0tWj.dm7YTc .i9lrp, .rFrNMe.k0tWj.dm7YTc .OabDMe { background-color: rgb(224, 96, 85); }

.whsOnd[disabled] { color: rgba(0, 0, 0, 0.38); }

.rFrNMe.dm7YTc .whsOnd[disabled] { color: rgba(255, 255, 255, 0.5); }

.whsOnd[disabled] ~ .i9lrp { background: none; border-bottom: 1px dotted rgba(0, 0, 0, 0.38); }

.OabDMe.Y2Zypf { animation: 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running quantumWizPaperInputRemoveUnderline; }

.rFrNMe.u3bW4e .OabDMe { animation: 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running quantumWizPaperInputAddUnderline; transform: scaleX(1); }

.rFrNMe.sdJrJc > .aCsJod { padding-top: 24px; }

.AxOyFc { transform-origin: left bottom; transition: color 0.3s cubic-bezier(0.4, 0, 0.2, 1) 0s, bottom, transform, -webkit-transform; color: rgba(0, 0, 0, 0.38); font: 400 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; pointer-events: none; position: absolute; bottom: 3px; left: 0px; width: 100%; }

.whsOnd:not([disabled]):focus ~ .AxOyFc, .whsOnd[badinput="true"] ~ .AxOyFc, .rFrNMe.CDELXb .AxOyFc, .rFrNMe.dLgj8b .AxOyFc { transform: scale(0.75) translateY(-39px); }

.whsOnd:not([disabled]):focus ~ .AxOyFc { color: rgb(51, 103, 214); }

.rFrNMe.dm7YTc .whsOnd:not([disabled]):focus ~ .AxOyFc { color: rgb(161, 194, 250); }

.rFrNMe.k0tWj .whsOnd:not([disabled]):focus ~ .AxOyFc { color: rgb(213, 0, 0); }

.ndJi5d { color: rgba(0, 0, 0, 0.38); font: 400 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; max-width: 100%; overflow: hidden; pointer-events: none; position: absolute; text-overflow: ellipsis; top: 2px; left: 0px; white-space: nowrap; }

.rFrNMe.CDELXb .ndJi5d { display: none; }

.K0Y8Se { -webkit-tap-highlight-color: transparent; font: 400 12px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 16px; margin-left: auto; padding-left: 16px; padding-top: 8px; pointer-events: none; opacity: 0.3; white-space: nowrap; }

.rFrNMe.dm7YTc .AxOyFc, .rFrNMe.dm7YTc .K0Y8Se, .rFrNMe.dm7YTc .ndJi5d { color: rgba(255, 255, 255, 0.7); }

.rFrNMe.Tyc9J { padding-bottom: 4px; }

.dEOOab, .ovnfwe:not(:empty) { -webkit-tap-highlight-color: transparent; -webkit-box-flex: 1; flex: 1 1 auto; font: 400 12px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; min-height: 16px; padding-top: 8px; }

.LXRPh { display: flex; }

.ovnfwe { pointer-events: none; }

.dEOOab { color: rgb(213, 0, 0); }

.rFrNMe.dm7YTc .dEOOab, .rFrNMe.dm7YTc.k0tWj .whsOnd:not([disabled]):focus ~ .AxOyFc { color: rgb(224, 96, 85); }

.ovnfwe { opacity: 0.3; }

.rFrNMe.dm7YTc .ovnfwe { color: rgba(255, 255, 255, 0.7); opacity: 1; }

.rFrNMe.k0tWj .ovnfwe, .rFrNMe:not(.k0tWj) .ovnfwe:not(:empty) + .dEOOab { display: none; }

@-webkit-keyframes quantumWizPaperInputRemoveUnderline { 
  0% { transform: scaleX(1); opacity: 1; }
  100% { transform: scaleX(1); opacity: 0; }
}

@keyframes quantumWizPaperInputRemoveUnderline { 
  0% { transform: scaleX(1); opacity: 1; }
  100% { transform: scaleX(1); opacity: 0; }
}

@-webkit-keyframes quantumWizPaperInputAddUnderline { 
  0% { transform: scaleX(0); }
  100% { transform: scaleX(1); }
}

@keyframes quantumWizPaperInputAddUnderline { 
  0% { transform: scaleX(0); }
  100% { transform: scaleX(1); }
}

.d1dlne, .Ax4B8 { display: flex; -webkit-box-flex: 1; flex: 1 1 0%; }

.L6J0Pc { -webkit-box-flex: 1; flex: 1 1 0%; }

.v5yLH, .v5yLH .d1dlne, .v5yLH .Ax4B8 { display: inline; }

.BBOA1c { position: absolute; height: 4px; bottom: 1px; left: 1px; right: 1px; overflow-x: hidden; background-color: rgb(255, 255, 255); display: none; }

.L6J0Pc.ge6pde .BBOA1c { display: block; }

.u3WVdc { position: absolute; right: 0px; left: 0px; z-index: 1; outline: none; overflow-y: auto; }

.u3WVdc[data-childcount="0"], .u3WVdc[data-expanded="false"] { display: none; }

.Cigftf { position: relative; top: -24px; }

.Ax4B8 { position: relative; }

.yNVtPc { position: absolute; left: 0px; width: 100%; opacity: 0.3; }

.Ax4B8, .yNVtPc { background-color: transparent; color: inherit; font: inherit; }

.d1dlne, .Ax4B8, .yNVtPc { height: 100%; }

.umNhxf { overflow-x: hidden; text-overflow: ellipsis; white-space: nowrap; }

.MkjOTb { cursor: default; }

.VOEIyf, .VOEIyf .jBmls, .oKubKe { font: 400 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(34, 34, 34); }

.VOEIyf { display: inline-block; height: 34px; line-height: 34px; }

.IjMZm { display: inline-block; height: auto; }

.VOEIyf .ZAGvjd { border-color: transparent; border-style: solid; border-width: 0px 1px; outline: none; }

.oKubKe, .VOEIyf .ZAGvjd { box-sizing: border-box; padding: 0px 16px; }

.VOEIyf .jBmls { box-sizing: border-box; padding: 8px 0px; border: 1px solid rgba(0, 0, 0, 0.2); background-color: rgb(255, 255, 255); border-radius: 0px 0px 2px 2px; box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; }

.oKubKe { line-height: 40px; }

.oKubKe[aria-selected="true"] { background-color: rgb(238, 238, 238); }

.oKubKe.RDPZE { color: rgba(0, 0, 0, 0.38); }

.SmXtye { margin: 7px 0px; border-top: 1px solid rgb(218, 218, 218); }

.D4D33b { overflow-x: hidden; text-overflow: ellipsis; white-space: nowrap; }

.oZ9DO { display: inline; }

.Pybrfb { fill: rgb(117, 117, 117); vertical-align: middle; }

.znqf0d { display: flex; line-height: 16px; padding-bottom: 8px; padding-top: 8px; }

.znqf0d .r3tIwf { -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; font-size: 16px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.znqf0d .r3tIwf .Ul51L { color: rgb(33, 33, 33); padding-top: 7px; }

.znqf0d .r3tIwf .VMD8Qc { color: rgb(117, 117, 117); padding-top: 3px; }

.znqf0d .RK4o7e { align-self: flex-end; -webkit-box-flex: 0; flex-grow: 0; flex-shrink: 0; height: 40px; padding: 4px 16px 4px 0px; }

.znqf0d .RhRPVd { height: 40px; width: 40px; border-radius: 50%; }

.RNHWXc .Pybrfb { margin-right: 16px; }

.pwHlAd { fill: rgb(255, 255, 255); height: 100%; vertical-align: middle; }

.DWfpSc, .ce4c1d { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; height: 34px; max-width: 100%; }

.DWn72e { height: 0px; overflow: hidden; visibility: hidden; }

.ce4c1d { position: relative; }

.Tfm4Hc .VOEIyf { height: 24px; line-height: 24px; max-width: 100%; }

.Tfm4Hc .oKubKe[aria-selected="true"] { outline: transparent solid 1px; }

.Tfm4Hc .d1dlne .ZAGvjd { -webkit-box-flex: 1; flex-grow: 1; padding: 0px; width: 0px; }

.Tfm4Hc .d1dlne[data-expanded="true"] .Ny5lGc { display: none; }

.Tfm4Hc .d1dlne .Ny5lGc { color: rgb(97, 97, 97); font-size: 14px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin-left: 1px; opacity: 1; pointer-events: none; width: calc(100% - 1px); z-index: 1; }

.Tfm4Hc .tWfTvb { bottom: 0px; left: 0px; position: absolute; width: 100%; }

.Tfm4Hc { max-width: 100%; }

.CjM6Fe { background-color: rgb(82, 100, 174); border-left: none; height: 36px; line-height: 34px; padding: 0px 4px; width: 36px; }

.CjM6Fe > .Pybrfb { vertical-align: middle; }

.mUbCce { user-select: none; transition: background 0.3s ease 0s; border: 0px; border-radius: 50%; cursor: pointer; display: inline-block; flex-shrink: 0; height: 48px; outline: none; overflow: hidden; position: relative; text-align: center; -webkit-tap-highlight-color: transparent; width: 48px; z-index: 0; }

.mUbCce > .TpQm9d { height: 48px; width: 48px; }

.mUbCce.u3bW4e, .mUbCce.qs41qe, .mUbCce.j7nIZb { transform: translateZ(0px); -webkit-mask-image: -webkit-radial-gradient(center, circle cover, white 100%, black 100%); }

.YYBxpf { border-radius: 0px; overflow: visible; }

.YYBxpf.u3bW4e, .YYBxpf.qs41qe, .YYBxpf.j7nIZb { -webkit-mask-image: none; }

.fKz7Od { color: rgba(0, 0, 0, 0.54); fill: rgba(0, 0, 0, 0.54); }

.p9Nwte { color: rgba(255, 255, 255, 0.75); fill: rgba(255, 255, 255, 0.75); }

.fKz7Od.u3bW4e { background-color: rgba(0, 0, 0, 0.12); }

.p9Nwte.u3bW4e { background-color: rgba(204, 204, 204, 0.25); }

.YYBxpf.u3bW4e { background-color: transparent; }

.VTBa7b { transform: translate(-50%, -50%) scale(0); transition: opacity 0.2s ease 0s, visibility 0s ease 0.2s, -webkit-transform 0s ease 0.2s; background-size: cover; left: 0px; opacity: 0; pointer-events: none; position: absolute; top: 0px; visibility: hidden; }

.YYBxpf.u3bW4e .VTBa7b { animation: 0.7s ease 0s infinite alternate none running quantumWizIconFocusPulse; height: 100%; left: 50%; top: 50%; width: 100%; visibility: visible; }

.mUbCce.qs41qe .VTBa7b { transform: translate(-50%, -50%) scale(2.2); opacity: 1; visibility: visible; }

.mUbCce.qs41qe.M9Bg4d .VTBa7b { transition: transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s, opacity 0.2s cubic-bezier(0, 0, 0.2, 1) 0s, -webkit-transform 0.3s cubic-bezier(0, 0, 0.2, 1) 0s; }

.mUbCce.j7nIZb .VTBa7b { transform: translate(-50%, -50%) scale(2.2); visibility: visible; }

.fKz7Od .VTBa7b { background-image: radial-gradient(circle farthest-side, rgba(0, 0, 0, 0.12), rgba(0, 0, 0, 0.12) 80%, rgba(0, 0, 0, 0) 100%); }

.p9Nwte .VTBa7b { background-image: radial-gradient(circle farthest-side, rgba(204, 204, 204, 0.25), rgba(204, 204, 204, 0.25) 80%, rgba(204, 204, 204, 0) 100%); }

.mUbCce.RDPZE { color: rgba(0, 0, 0, 0.26); fill: rgba(0, 0, 0, 0.26); cursor: default; }

.p9Nwte.RDPZE { color: rgba(255, 255, 255, 0.5); fill: rgba(255, 255, 255, 0.5); }

.xjKiLb { position: relative; top: 50%; }

.xjKiLb > span { display: inline-block; position: relative; }

.SPwuPd { -webkit-box-align: center; align-items: center; display: flex; height: 24px; margin-bottom: 3px; margin-right: 3px; overflow: hidden; padding-left: 2px; white-space: nowrap; position: relative; z-index: 1; }

.tRMgEc { border-radius: 50%; -webkit-user-drag: none; }

.HYyewd { color: rgb(97, 97, 97); font: 500 12px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin-left: 8px; overflow-x: hidden; text-overflow: ellipsis; }

.WqfY4c { height: 32px; width: 32px; }

.SPwuPd.cTDLLd { background: rgb(255, 255, 255); border: 1px solid rgb(224, 224, 224); border-radius: 16px; }

.SPwuPd.o1yOod { background: rgb(245, 245, 245); border: 1px solid rgb(250, 218, 128); border-radius: 3px; }

.SPwuPd.ui9xvd > .HYyewd { border-bottom: 2px dotted rgb(211, 47, 47); }

.Tezzlf > .HYyewd { margin-right: 8px; }

.Cbzx4b { -webkit-box-align: center; align-items: center; border-radius: 50%; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; font: 400 13px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 20px; -webkit-box-pack: center; justify-content: center; opacity: 0.6; text-transform: uppercase; width: 20px; }

.mElJdc { fill: rgb(229, 57, 53); padding-left: 1px; }

.FKF6mc, .FKF6mc:focus { display: block; outline: none; text-decoration: none; }

.FKF6mc:visited { fill: inherit; stroke: inherit; }

.U26fgb.u3bW4e { outline: transparent solid 1px; }

.w6DEz { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-flex: 1; flex: 1 1 auto; flex-wrap: wrap; -webkit-box-pack: start; justify-content: flex-start; max-height: 100%; min-height: 24px; overflow: hidden auto; width: 100%; }

.IHB8eb { -webkit-box-align: center; align-items: center; display: inline-flex; -webkit-box-flex: 0; flex: 0 0 auto; flex-wrap: wrap; -webkit-box-pack: start; justify-content: flex-start; max-height: 100%; max-width: 100%; min-height: 24px; overflow-y: auto; width: 100%; }

.IHB8eb .u3WVdc { z-index: 2000; }

.ARQdkc, .ZeowYe { -webkit-box-flex: 1; flex-grow: 1; padding-bottom: 0px; }

.ARQdkc { cursor: text; display: flex; -webkit-box-pack: justify; justify-content: space-between; max-width: 100%; position: relative; }

.qH6atb, .eONaNc { display: block; -webkit-box-flex: 0; flex: 0 0 auto; }

.ARQdkc.DHpaLb .ZeowYe { display: none; }

.zVw2Qe { box-sizing: border-box; display: none; -webkit-box-flex: 1; flex: 1 1 auto; height: 34px; line-height: 34px; width: 0px; }

.ARQdkc.DHpaLb .zVw2Qe { display: inline-flex; }

.R7dqcc { background-color: transparent; border: none; color: inherit; font: inherit; height: 100%; outline: none; padding: 0px; width: 100%; }

.ARQdkc .ZAGvjd { border: none; }

.QsGMEc { background-color: rgb(255, 255, 255); border-radius: 0px 0px 2px 2px; border: 1px solid rgba(0, 0, 0, 0.2); box-shadow: rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px, rgba(0, 0, 0, 0.2) 0px 5px 5px -3px; box-sizing: border-box; display: none; left: 0px; padding: 8px 0px; position: absolute; right: 0px; top: 100%; z-index: 0; }

.zVw2Qe.KrQ13 .QsGMEc { display: block; z-index: 1; }

.r5czLc { line-height: 24px; overflow: hidden; padding-left: 16px; white-space: normal; }

.GGoold { -webkit-box-align: center; align-items: center; display: flex; }

.r5czLc.r5czLc { color: rgb(128, 134, 139); }

.itOdAb { fill: rgb(128, 134, 139); }

.tFoQfe { background: canvas; border: 1px solid transparent; border-radius: 8px; box-sizing: border-box; display: block; max-height: 100%; max-width: 100%; pointer-events: auto; z-index: 0; }

.tFoQfe:focus { outline: none; }

.tFoQfe:focus-visible { outline: initial; }

.Q5UMwc { display: block; height: 100%; left: 0px; pointer-events: auto; position: fixed; top: 0px; width: 100%; z-index: 0; }

.PPAvie { -webkit-box-align: center; align-items: center; inset: 0px; display: flex; -webkit-box-pack: center; justify-content: center; pointer-events: none; position: absolute; z-index: 0; }

.Ae8Td { animation: 0.15s linear 0s 1 normal backwards running drive-elements-dialog-fade-in; background: var(--dt-scrim,rgba(32,33,36,.6)); }

[hidden] .Ae8Td { animation: 75ms linear 0s 1 normal both running drive-elements-dialog-fade-out; }

.iYu4xd { background: var(--dt-surface3,#fff); border: 1px solid transparent; border-radius: 8px; box-shadow: var(--dt-surface3-shadow,0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15)); box-sizing: border-box; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; margin: 24px; max-width: 512px; min-width: 320px; padding-top: 24px; pointer-events: auto; position: relative; transform-origin: center center; z-index: 1; }

.vhoiae .iYu4xd { background: var(--dt-background,#fff); }

@media screen and (max-width: 320px) {
  .iYu4xd { margin: 12px; max-width: 100%; min-width: 0px; }
}

.iYu4xd { animation: 75ms linear 0s 1 normal backwards running drive-elements-dialog-fade-in, 0.15s cubic-bezier(0, 0, 0.2, 1) 0s 1 normal backwards running drive-elements-dialog-transform; }

.iYu4xd.yoBxB { max-width: 832px; padding-top: 0px; }

[hidden] .iYu4xd { animation: 75ms linear 0s 1 normal forwards running drive-elements-dialog-fade-out; }

.ROcXFc { box-sizing: border-box; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; max-height: 100%; min-height: 0px; width: 100%; }

.FidVJb { box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); cursor: default; -webkit-box-flex: 0; flex: 0 0 auto; font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 1.375rem; font-weight: 500; line-height: 1.5rem; margin-bottom: 12px; margin-top: 0px; padding: 0px 24px; }

.vhoiae .FidVJb, .X9XeLb .FidVJb, .cWKK1c .FidVJb, .aJfoSc .FidVJb, .TOb6Ze .FidVJb { font: var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-headline-small-spacing,0); margin-bottom: 16px; }

.FidVJb.cd29Sd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; text-align: center; }

.kOD2fb { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); cursor: default; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 auto; margin-bottom: 12px; overflow: auto; padding: 0px; width: 100%; }

.OsLnq { box-sizing: border-box; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-pack: end; justify-content: flex-end; padding: 8px 16px 8px 0px; }

.OsLnq.IRlIld { padding: 8px 24px 16px 0px; }

.uAkPhe.vKmmhc, .wnagdd.vKmmhc, .oB1s2d.vKmmhc { margin-left: 8px; }

.ThEHqd { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-pack: center; justify-content: center; }

.zsVT8c { color: var(--dt-on-surface,rgb(60,64,67)); fill: currentcolor; font-size: 24px; margin-bottom: 12px; }

.zsVT8c.kphldf { color: var(--dt-error,rgb(217,48,37)); }

.zsVT8c.sj692e { color: var(--dt-primary,rgb(26,115,232)); }

.zsVT8c.IY5c4e { color: var(--dt-tertiary,rgb(24,128,56)); }

.zsVT8c.rNe0id { color: var(--dt-warning,rgb(249,171,0)); }

.ELTUEc { color: var(--dt-on-surface,rgb(60,64,67)); display: flex; fill: currentcolor; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; font-size: 1.5rem; -webkit-box-pack: center; justify-content: center; margin-bottom: 0.75rem; }

.ELTUEc.kphldf { color: var(--dt-error,rgb(217,48,37)); }

.ELTUEc.sj692e { color: var(--dt-primary,rgb(26,115,232)); }

.ELTUEc.IY5c4e { color: var(--dt-tertiary,rgb(24,128,56)); }

.ELTUEc.rNe0id { color: var(--dt-warning,rgb(249,171,0)); }

.jOirTd { -webkit-box-flex: 0; flex: 0 0 auto; }

.P6NGpd { color: var(--dt-primary-container-link,rgb(25,103,210)); }

.BvVDgb { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); background: var(--dt-surface-variant,rgb(241,243,244)); border-bottom: 1px solid var(--dt-outline,rgb(128,134,139)); border-left: 1px solid var(--dt-outline,rgb(128,134,139)); border-radius: 0px 6px 0px 0px; box-sizing: border-box; color: var(--dt-on-surface,rgb(60,64,67)); cursor: default; max-width: 320px; padding: 1.5rem 1.5rem 0.75rem; }

.U5qczb { display: flex; }

.HY9Yxe { -webkit-box-flex: 1; flex: 1 1 auto; }

.HY9Yxe.yoBxB { padding-top: 24px; }

.y42Lxf { position: absolute; top: 0px; right: 0px; }

@-webkit-keyframes drive-elements-dialog-fade-in { 
  0% { opacity: 0; }
  100% { opacity: 1; }
}

@keyframes drive-elements-dialog-fade-in { 
  0% { opacity: 0; }
  100% { opacity: 1; }
}

@-webkit-keyframes drive-elements-dialog-fade-out { 
  0% { opacity: 1; visibility: visible; }
  99.998% { opacity: 0; visibility: visible; }
  99.999%, 100% { opacity: 0; visibility: hidden; }
}

@keyframes drive-elements-dialog-fade-out { 
  0% { opacity: 1; visibility: visible; }
  99.998% { opacity: 0; visibility: visible; }
  99.999%, 100% { opacity: 0; visibility: hidden; }
}

@-webkit-keyframes drive-elements-dialog-transform { 
  0% { transform: none; }
  1% { transform: scale(0.8); }
  100% { transform: scale(1); }
}

@keyframes drive-elements-dialog-transform { 
  0% { transform: none; }
  1% { transform: scale(0.8); }
  100% { transform: scale(1); }
}

.FlWAte { width: 600px; max-width: 600px; height: 550px; padding-top: 12px; }

.HnJMoe { box-sizing: border-box; display: flex; flex-direction: row; height: 460px; padding-right: 8px; width: 100%; }

.axuJCe { flex: 0 0 220px; overflow: hidden auto; }

.HnJMoe.EBwNne .axuJCe { display: none; }

.EEauGd { margin-left: 8px; flex: 1 1 60%; position: relative; overflow-y: auto; }

.IIpXyc { border-radius: 0px 35px 35px 0px; box-sizing: border-box; display: flex; margin-top: 8px; overflow-x: hidden; width: 100%; padding: 4px 16px 4px 22px; }

.IIpXyc.Er3Sgf { border: 1px solid transparent; background: var(--dt-primary-container,#e8f0fe); }

.IIpXyc.UQXU5c { color: var(--dt-on-surface,#3c4043); opacity: 0.38; }

.uDfb0b { margin-top: 8px; }

.nYTocd { margin-bottom: -12px; }

.nRg5rb { display: flex; align-items: center; }

.pBhHJc { margin-left: auto; margin-right: -12px; }

.pBhHJc:focus::before, .pBhHJc:hover::before { border: 1px dashed transparent; border-radius: 50%; inset: 0px; content: ""; margin: 1px; position: absolute; }

.I8jRHe { fill: var(--dt-background,#fff); margin-right: 1px; }

.jJrJwd { align-items: center; background: var(--dt-primary-action-state-layer,#1967d2); border-radius: 50%; display: flex; height: 28px; justify-content: center; margin-right: 5px; width: 28px; }

.qBWx0d { overflow-x: hidden; }

.t3R3ld { overflow-x: hidden; text-overflow: ellipsis; white-space: nowrap; }

.x1qPs { height: 16px; padding: 2px 8px 0px 0px; }

.oT1Ike { width: 16px; }

.ycrW9 { align-content: center; -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; list-style: none; margin: 0px; max-height: 100%; max-width: 100%; padding: 0px; }

.ycrW9:focus { outline: none; }

.ycrW9[aria-orientation="horizontal"] { -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.BmS7Jf { }

.BmS7Jf:hover, .BmS7Jf:active, .BmS7Jf:focus-within { }

.BmS7Jf::-webkit-scrollbar { background-color: transparent; border-radius: 0px; height: 8px; width: 8px; }

.BmS7Jf::-webkit-scrollbar-thumb { background-color: transparent; }

.BmS7Jf::-webkit-scrollbar-thumb:active { background-color: transparent; }

.BmS7Jf:hover::-webkit-scrollbar { background-color: transparent; }

.BmS7Jf:hover::-webkit-scrollbar-thumb, .BmS7Jf:focus-within::-webkit-scrollbar-thumb { background-color: rgba(95, 99, 104, 0.2); background-clip: padding-box; border-radius: 0px; padding: 100px 0px 0px; }

@media (forced-colors: active) {
  .BmS7Jf:hover::-webkit-scrollbar-thumb, .BmS7Jf:focus-within::-webkit-scrollbar-thumb { background-color: canvastext; }
}

.BmS7Jf::-webkit-scrollbar-thumb:hover { background-color: rgba(95, 99, 104, 0.2); }

@media (forced-colors: active) {
  .BmS7Jf::-webkit-scrollbar-thumb:hover { background-color: canvastext; }
}

@media (forced-colors: active) {
}

.BmS7Jf::-webkit-scrollbar-corner { background: transparent; }

.gKD1Qc::-webkit-scrollbar { width: 12px; }

.gKD1Qc::-webkit-scrollbar-button { height: 0px; width: 0px; }

.gKD1Qc::-webkit-scrollbar-thumb, .gKD1Qc::-webkit-scrollbar-thumb:hover, .gKD1Qc::-webkit-scrollbar-thumb:active { background-color: rgba(66, 133, 244, 0.32); }

@media (forced-colors: active) {
  .gKD1Qc::-webkit-scrollbar-thumb, .gKD1Qc::-webkit-scrollbar-thumb:hover, .gKD1Qc::-webkit-scrollbar-thumb:active { background-color: canvastext; }
}

.gKD1Qc.hpDt6e::-webkit-scrollbar-thumb { border-radius: 4px; }

.gKD1Qc.kbeFSb::-webkit-scrollbar-thumb { border-radius: 4px 0px 0px 4px; }

.ZACE2c { -webkit-box-align: center; align-items: center; inset: 0px; display: flex; height: 100%; -webkit-box-pack: center; justify-content: center; pointer-events: none; position: fixed; width: 100%; z-index: 2300; }

.ZACE2c:not(.eO2Zfd) { display: none; }

.mC2T2 { inset: 0px; display: block; pointer-events: none; position: absolute; visibility: hidden; z-index: 0; }

.xmQMab { pointer-events: auto; z-index: 1; }

.VfPpkd-MPu53c { padding: calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2); margin: calc((var(--mdc-checkbox-touch-target-size, 40px) - 40px)/2); }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c .VfPpkd-OYHm6b::after { background-color: var(--mdc-ripple-color,#000); }

.VfPpkd-MPu53c:hover .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786)); }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:hover .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786)); }

.VfPpkd-MPu53c .VfPpkd-YQoJzd { top: calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2); left: calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe { top: calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2); right: calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2); left: calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2); width: var(--mdc-checkbox-touch-target-size,40px); height: var(--mdc-checkbox-touch-target-size,40px); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54)); background-color: transparent; }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); background-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); }

@-webkit-keyframes mdc-checkbox-fade-in-background-8A000000FF01878600000000FF018786 { 
  0% { border-color: var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54)); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); background-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); }
}

@keyframes mdc-checkbox-fade-in-background-8A000000FF01878600000000FF018786 { 
  0% { border-color: var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54)); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); background-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); }
}

@-webkit-keyframes mdc-checkbox-fade-out-background-8A000000FF01878600000000FF018786 { 
  0%, 80% { border-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); background-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); }
  100% { border-color: var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54)); background-color: transparent; }
}

@keyframes mdc-checkbox-fade-out-background-8A000000FF01878600000000FF018786 { 
  0%, 80% { border-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); background-color: var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786)); }
  100% { border-color: var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54)); background-color: transparent; }
}

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-in-background-8A000000FF01878600000000FF018786; }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-out-background-8A000000FF01878600000000FF018786; }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-disabled-color,rgba(0,0,0,.38)); background-color: transparent; }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:checked ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"][disabled] ~ .VfPpkd-YQoJzd { border-color: transparent; background-color: var(--mdc-checkbox-disabled-color,rgba(0,0,0,.38)); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-ink-color,#fff); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-ink-color,#fff); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-ink-color,#fff); }

.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-ink-color,#fff); }

@-webkit-keyframes mdc-checkbox-unchecked-checked-checkmark-path { 
  0%, 50% { stroke-dashoffset: 29.7833; }
  50% { animation-timing-function: cubic-bezier(0, 0, 0.2, 1); }
  100% { stroke-dashoffset: 0; }
}

@keyframes mdc-checkbox-unchecked-checked-checkmark-path { 
  0%, 50% { stroke-dashoffset: 29.7833; }
  50% { animation-timing-function: cubic-bezier(0, 0, 0.2, 1); }
  100% { stroke-dashoffset: 0; }
}

@-webkit-keyframes mdc-checkbox-unchecked-indeterminate-mixedmark { 
  0%, 68.2% { transform: scaleX(0); }
  68.2% { animation-timing-function: cubic-bezier(0, 0, 0, 1); }
  100% { transform: scaleX(1); }
}

@keyframes mdc-checkbox-unchecked-indeterminate-mixedmark { 
  0%, 68.2% { transform: scaleX(0); }
  68.2% { animation-timing-function: cubic-bezier(0, 0, 0, 1); }
  100% { transform: scaleX(1); }
}

@-webkit-keyframes mdc-checkbox-checked-unchecked-checkmark-path { 
  0% { animation-timing-function: cubic-bezier(0.4, 0, 1, 1); opacity: 1; stroke-dashoffset: 0; }
  100% { opacity: 0; stroke-dashoffset: -29.7833; }
}

@keyframes mdc-checkbox-checked-unchecked-checkmark-path { 
  0% { animation-timing-function: cubic-bezier(0.4, 0, 1, 1); opacity: 1; stroke-dashoffset: 0; }
  100% { opacity: 0; stroke-dashoffset: -29.7833; }
}

@-webkit-keyframes mdc-checkbox-checked-indeterminate-checkmark { 
  0% { animation-timing-function: cubic-bezier(0, 0, 0.2, 1); transform: rotate(0deg); opacity: 1; }
  100% { transform: rotate(45deg); opacity: 0; }
}

@keyframes mdc-checkbox-checked-indeterminate-checkmark { 
  0% { animation-timing-function: cubic-bezier(0, 0, 0.2, 1); transform: rotate(0deg); opacity: 1; }
  100% { transform: rotate(45deg); opacity: 0; }
}

@-webkit-keyframes mdc-checkbox-indeterminate-checked-checkmark { 
  0% { animation-timing-function: cubic-bezier(0.14, 0, 0, 1); transform: rotate(45deg); opacity: 0; }
  100% { transform: rotate(1turn); opacity: 1; }
}

@keyframes mdc-checkbox-indeterminate-checked-checkmark { 
  0% { animation-timing-function: cubic-bezier(0.14, 0, 0, 1); transform: rotate(45deg); opacity: 0; }
  100% { transform: rotate(1turn); opacity: 1; }
}

@-webkit-keyframes mdc-checkbox-checked-indeterminate-mixedmark { 
  0% { transform: rotate(-45deg); opacity: 0; }
  100% { transform: rotate(0deg); opacity: 1; }
}

@keyframes mdc-checkbox-checked-indeterminate-mixedmark { 
  0% { transform: rotate(-45deg); opacity: 0; }
  100% { transform: rotate(0deg); opacity: 1; }
}

@-webkit-keyframes mdc-checkbox-indeterminate-checked-mixedmark { 
  0% { animation-timing-function: cubic-bezier(0.14, 0, 0, 1); transform: rotate(0deg); opacity: 1; }
  100% { transform: rotate(315deg); opacity: 0; }
}

@keyframes mdc-checkbox-indeterminate-checked-mixedmark { 
  0% { animation-timing-function: cubic-bezier(0.14, 0, 0, 1); transform: rotate(0deg); opacity: 1; }
  100% { transform: rotate(315deg); opacity: 0; }
}

@-webkit-keyframes mdc-checkbox-indeterminate-unchecked-mixedmark { 
  0% { animation-timing-function: linear; transform: scaleX(1); opacity: 1; }
  32.8%, 100% { transform: scaleX(0); opacity: 0; }
}

@keyframes mdc-checkbox-indeterminate-unchecked-mixedmark { 
  0% { animation-timing-function: linear; transform: scaleX(1); opacity: 1; }
  32.8%, 100% { transform: scaleX(0); opacity: 0; }
}

.VfPpkd-MPu53c { display: inline-block; position: relative; -webkit-box-flex: 0; flex: 0 0 18px; box-sizing: content-box; width: 18px; height: 18px; line-height: 0; white-space: nowrap; cursor: pointer; vertical-align: bottom; }

.VfPpkd-MPu53c[hidden] { display: none; }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec, .VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec { pointer-events: none; border: 2px solid transparent; border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: 100%; width: 100%; }

@media screen and (forced-colors: active) {
  .VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec, .VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec { border-color: canvastext; }
}

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec::after, .VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec::after { content: ""; border: 2px solid transparent; border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec::after, .VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec::after { border-color: canvastext; }
}

@media (-ms-high-contrast:none) {
  .VfPpkd-MPu53c .VfPpkd-sMek6-LhBDec { display: none; }
}

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .VfPpkd-SJnn3d { margin: 0px 1px; }
}

.VfPpkd-MPu53c-OWXEXe-OWB6Me { cursor: default; pointer-events: none; }

.VfPpkd-YQoJzd { display: inline-flex; position: absolute; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; box-sizing: border-box; width: 18px; height: 18px; border: 2px solid currentcolor; border-radius: 2px; background-color: transparent; pointer-events: none; will-change: background-color, border-color; transition: background-color 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms, border-color 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-HUofsb { position: absolute; inset: 0px; width: 100%; opacity: 0; transition: opacity 0.18s cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb { opacity: 1; }

.VfPpkd-HUofsb-Jt5cK { transition: stroke-dashoffset 0.18s cubic-bezier(0.4, 0, 0.6, 1) 0ms; stroke: currentcolor; stroke-width: 3.12px; stroke-dashoffset: 29.7833; stroke-dasharray: 29.7833; }

.VfPpkd-SJnn3d { width: 100%; height: 0px; transform: scaleX(0) rotate(0deg); border-width: 1px; border-style: solid; opacity: 0; transition: opacity 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms, transform 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms, -webkit-transform 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-YQoJzd, .VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-YQoJzd, .VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-YQoJzd, .VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-YQoJzd { animation-duration: 0.18s; animation-timing-function: linear; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-HUofsb-Jt5cK { animation: 0.18s linear 0s 1 normal none running mdc-checkbox-unchecked-checked-checkmark-path; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-SJnn3d { animation: 90ms linear 0s 1 normal none running mdc-checkbox-unchecked-indeterminate-mixedmark; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-HUofsb-Jt5cK { animation: 90ms linear 0s 1 normal none running mdc-checkbox-checked-unchecked-checkmark-path; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-A9y3zc .VfPpkd-HUofsb { animation: 90ms linear 0s 1 normal none running mdc-checkbox-checked-indeterminate-checkmark; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-A9y3zc .VfPpkd-SJnn3d { animation: 90ms linear 0s 1 normal none running mdc-checkbox-checked-indeterminate-mixedmark; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-barxie .VfPpkd-HUofsb { animation: 0.5s linear 0s 1 normal none running mdc-checkbox-indeterminate-checked-checkmark; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-barxie .VfPpkd-SJnn3d { animation: 0.5s linear 0s 1 normal none running mdc-checkbox-indeterminate-checked-mixedmark; transition: none 0s ease 0s; }

.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-SJnn3d { animation: 0.3s linear 0s 1 normal none running mdc-checkbox-indeterminate-unchecked-mixedmark; transition: none 0s ease 0s; }

.VfPpkd-muHVFf-bMcfAe:checked ~ .VfPpkd-YQoJzd, .VfPpkd-muHVFf-bMcfAe:indeterminate ~ .VfPpkd-YQoJzd, .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"] ~ .VfPpkd-YQoJzd { transition: border-color 90ms cubic-bezier(0, 0, 0.2, 1) 0ms, background-color 90ms cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-muHVFf-bMcfAe:checked ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK, .VfPpkd-muHVFf-bMcfAe:indeterminate ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK, .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"] ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK { stroke-dashoffset: 0; }

.VfPpkd-muHVFf-bMcfAe { position: absolute; margin: 0px; padding: 0px; opacity: 0; cursor: inherit; }

.VfPpkd-muHVFf-bMcfAe:disabled { cursor: default; pointer-events: none; }

.VfPpkd-MPu53c-OWXEXe-dgl2Hf { margin: calc((var(--mdc-checkbox-state-layer-size, 48px) - var(--mdc-checkbox-state-layer-size, 40px))/2); }

.VfPpkd-MPu53c-OWXEXe-dgl2Hf .VfPpkd-muHVFf-bMcfAe { top: calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2); right: calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2); left: calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2); width: var(--mdc-checkbox-state-layer-size,48px); height: var(--mdc-checkbox-state-layer-size,48px); }

.VfPpkd-muHVFf-bMcfAe:checked ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { transition: opacity 0.18s cubic-bezier(0, 0, 0.2, 1) 0ms, transform 0.18s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.18s cubic-bezier(0, 0, 0.2, 1) 0ms; opacity: 1; }

.VfPpkd-muHVFf-bMcfAe:checked ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { transform: scaleX(1) rotate(-45deg); }

.VfPpkd-muHVFf-bMcfAe:indeterminate ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb, .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"] ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { transform: rotate(45deg); opacity: 0; transition: opacity 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms, transform 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms, -webkit-transform 90ms cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-muHVFf-bMcfAe:indeterminate ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d, .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"] ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { transform: scaleX(1) rotate(0deg); opacity: 1; }

.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-YQoJzd, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb-Jt5cK, .VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-SJnn3d { transition: none 0s ease 0s; }

.VfPpkd-MPu53c { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c .VfPpkd-OYHm6b::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-OYHm6b::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-OYHm6b::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-OYHm6b::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c .VfPpkd-OYHm6b::after { top: 0px; left: 0px; width: 100%; height: 100%; }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-MPu53c { z-index: 0; }

.VfPpkd-MPu53c .VfPpkd-OYHm6b::before, .VfPpkd-MPu53c .VfPpkd-OYHm6b::after { z-index: var(--mdc-ripple-z-index,-1); }

.VfPpkd-OYHm6b { position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; pointer-events: none; }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-disabled-unselected-icon-color,GrayText); background-color: transparent; }
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:checked ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate ~ .VfPpkd-YQoJzd, .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"][disabled] ~ .VfPpkd-YQoJzd { border-color: graytext; background-color: var(--mdc-checkbox-disabled-selected-icon-color,GrayText); }
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-selected-checkmark-color,ButtonText); }
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-selected-checkmark-color,ButtonText); }
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace); }
  .VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace); }
}

.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-disabled-unselected-icon-color,rgba(60,64,67,.38)); background-color: transparent; }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:checked ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"][disabled] ~ .VfPpkd-YQoJzd { border-color: transparent; background-color: var(--mdc-checkbox-disabled-selected-icon-color,rgba(60,64,67,.38)); }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-selected-checkmark-color,#fff); }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-selected-checkmark-color,#fff); }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-disabled-selected-checkmark-color,#fff); }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-disabled-selected-checkmark-color,#fff); }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-unselected-icon-color,#5f6368); background-color: transparent; }

.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); background-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); }

@-webkit-keyframes mdc-checkbox-fade-in-background-FF5F6368FF1A73E800000000FF1A73E8 { 
  0% { border-color: var(--mdc-checkbox-unselected-icon-color,#5f6368); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); background-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); }
}

@keyframes mdc-checkbox-fade-in-background-FF5F6368FF1A73E800000000FF1A73E8 { 
  0% { border-color: var(--mdc-checkbox-unselected-icon-color,#5f6368); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); background-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); }
}

@-webkit-keyframes mdc-checkbox-fade-out-background-FF5F6368FF1A73E800000000FF1A73E8 { 
  0%, 80% { border-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); background-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); }
  100% { border-color: var(--mdc-checkbox-unselected-icon-color,#5f6368); background-color: transparent; }
}

@keyframes mdc-checkbox-fade-out-background-FF5F6368FF1A73E800000000FF1A73E8 { 
  0%, 80% { border-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); background-color: var(--mdc-checkbox-selected-icon-color,#1a73e8); }
  100% { border-color: var(--mdc-checkbox-unselected-icon-color,#5f6368); background-color: transparent; }
}

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-in-background-FF5F6368FF1A73E800000000FF1A73E8; }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-out-background-FF5F6368FF1A73E800000000FF1A73E8; }

.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-unselected-hover-icon-color,#202124); background-color: transparent; }

.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); }

@-webkit-keyframes mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6 { 
  0% { border-color: var(--mdc-checkbox-unselected-hover-icon-color,#202124); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); }
}

@-webkit-keyframes mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6 { 
  0%, 80% { border-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-hover-icon-color,#174ea6); }
  100% { border-color: var(--mdc-checkbox-unselected-hover-icon-color,#202124); background-color: transparent; }
}

.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-unselected-focus-icon-color,#202124); background-color: transparent; }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-selected-focus-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-focus-icon-color,#174ea6); }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-unselected-pressed-icon-color,#202124); background-color: transparent; }

.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked ~ .VfPpkd-YQoJzd, .Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"]:enabled ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); }

@keyframes mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6 { 
  0% { border-color: var(--mdc-checkbox-unselected-pressed-icon-color,#202124); background-color: transparent; }
  50% { border-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); }
}

@keyframes mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6 { 
  0%, 80% { border-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); background-color: var(--mdc-checkbox-selected-pressed-icon-color,#174ea6); }
  100% { border-color: var(--mdc-checkbox-unselected-pressed-icon-color,#202124); background-color: transparent; }
}

.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd, .Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd { animation-name: mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6; }

.Ne8lhe .VfPpkd-OYHm6b::before, .Ne8lhe .VfPpkd-OYHm6b::after { background-color: var(--mdc-checkbox-unselected-hover-state-layer-color,#3c4043); }

.Ne8lhe:hover .VfPpkd-OYHm6b::before, .Ne8lhe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before { opacity: var(--mdc-checkbox-unselected-hover-state-layer-opacity,.04); }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before, .Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before { transition-duration: 75ms; opacity: var(--mdc-checkbox-unselected-focus-state-layer-opacity,.12); }

.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after { transition: opacity 0.15s linear 0s; }

.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after { transition-duration: 75ms; opacity: var(--mdc-checkbox-unselected-pressed-state-layer-opacity,.1); }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-checkbox-unselected-pressed-state-layer-opacity,0.1); }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before, .Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after { background-color: var(--mdc-checkbox-selected-hover-state-layer-color,#1a73e8); }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:hover .VfPpkd-OYHm6b::before, .Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before { opacity: var(--mdc-checkbox-selected-hover-state-layer-opacity,.04); }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before, .Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before { transition-duration: 75ms; opacity: var(--mdc-checkbox-selected-focus-state-layer-opacity,.12); }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after { transition: opacity 0.15s linear 0s; }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after { transition-duration: 75ms; opacity: var(--mdc-checkbox-selected-pressed-state-layer-opacity,.1); }

.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-checkbox-selected-pressed-state-layer-opacity,0.1); }

.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before, .Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after { background-color: var(--mdc-checkbox-selected-hover-state-layer-color,#1a73e8); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate="true"]) ~ .VfPpkd-YQoJzd { border-color: var(--mdc-checkbox-disabled-unselected-icon-color,GrayText); background-color: transparent; }
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:checked ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate ~ .VfPpkd-YQoJzd, .Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate="true"][disabled] ~ .VfPpkd-YQoJzd { border-color: graytext; background-color: var(--mdc-checkbox-disabled-selected-icon-color,GrayText); }
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-selected-checkmark-color,ButtonText); }
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-selected-checkmark-color,ButtonText); }
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-HUofsb { color: var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace); }
  .Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled ~ .VfPpkd-YQoJzd .VfPpkd-SJnn3d { border-color: var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace); }
}

.az2ine { will-change: unset; }

.VfPpkd-I9GLp-yrriRe { display: inline-flex; -webkit-box-align: center; align-items: center; vertical-align: middle; }

.VfPpkd-I9GLp-yrriRe[hidden] { display: none; }

.VfPpkd-I9GLp-yrriRe > label { margin-left: 0px; margin-right: auto; padding-left: 4px; padding-right: 0px; -webkit-box-ordinal-group: 1; order: 0; }

[dir="rtl"] .VfPpkd-I9GLp-yrriRe > label, .VfPpkd-I9GLp-yrriRe > label[dir="rtl"] { margin-left: auto; margin-right: 0px; }

[dir="rtl"] .VfPpkd-I9GLp-yrriRe > label, .VfPpkd-I9GLp-yrriRe > label[dir="rtl"] { padding-left: 0px; padding-right: 4px; }

.VfPpkd-I9GLp-yrriRe-OWXEXe-WrakWd > label { text-overflow: ellipsis; overflow: hidden; white-space: nowrap; }

.VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d > label { margin-left: auto; margin-right: 0px; padding-left: 0px; padding-right: 4px; order: -1; }

[dir="rtl"] .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d > label, .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d > label[dir="rtl"] { margin-left: 0px; margin-right: auto; }

[dir="rtl"] .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d > label, .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d > label[dir="rtl"] { padding-left: 4px; padding-right: 0px; }

.VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL { -webkit-box-pack: justify; justify-content: space-between; }

.VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL > label { margin: 0px; }

[dir="rtl"] .VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL > label, .VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL > label[dir="rtl"] { margin: 0px; }

.VfPpkd-I9GLp-yrriRe { font-family: var(--mdc-form-field-label-text-font,Roboto,sans-serif); line-height: var(--mdc-form-field-label-text-line-height,1.25rem); font-size: var(--mdc-form-field-label-text-size,.875rem); font-weight: var(--mdc-form-field-label-text-weight,400); letter-spacing: var(--mdc-form-field-label-text-tracking,.0178571429em); color: var(--mdc-form-field-label-text-color,var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))); }

.MlG5Jc { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; }

.MlG5Jc gm-checkbox[disabled] ~ .VfPpkd-V67aGc, .MlG5Jc gm-radio[disabled] ~ .VfPpkd-V67aGc, .MlG5Jc .VfPpkd-MPu53c-OWXEXe-OWB6Me ~ .VfPpkd-V67aGc, .MlG5Jc .VfPpkd-GCYh9b-OWXEXe-OWB6Me ~ .VfPpkd-V67aGc { color: rgb(95, 99, 104); }

.p9IRvd { box-sizing: border-box; max-height: 100%; max-width: 100%; padding: 0px 1.5rem; white-space: pre-line; }

.Q7xaL { left: -1rem; margin-top: 0.5rem; position: relative; }

.Q7xaL .VfPpkd-muHVFf-bMcfAe:focus ~ .VfPpkd-OYHm6b { outline: transparent solid 1px; }

.fsrxTe { box-sizing: border-box; max-height: 100%; max-width: 100%; padding: 0px 1.5rem; white-space: pre-line; }

.UGmH4e { box-sizing: border-box; max-height: 100%; max-width: 100%; padding: 0.25rem 1.25rem 0px; }

.Mh0NNb { background-color: rgb(50, 50, 50); bottom: 0px; box-sizing: border-box; box-shadow: rgba(0, 0, 0, 0.14) 0px 6px 10px 0px, rgba(0, 0, 0, 0.12) 0px 1px 18px 0px, rgba(0, 0, 0, 0.2) 0px 3px 5px -1px; color: rgb(255, 255, 255); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; font-size: 14px; left: 0px; min-height: 48px; position: fixed; right: 0px; transform: translate(0px, 100%); visibility: hidden; z-index: 99999; }

.M6tHv { -webkit-box-align: center; align-items: center; align-content: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; min-height: inherit; padding: 0px; }

.aGJE1b { -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; line-height: normal; overflow: hidden; padding: 14px 24px; text-overflow: ellipsis; word-break: break-word; }

.x95qze { align-self: center; color: rgb(238, 255, 65); -webkit-box-flex: 0; flex-grow: 0; flex-shrink: 0; float: right; text-transform: uppercase; font-weight: 500; display: inline-block; cursor: pointer; outline: none; padding: 14px 24px; }

.KYZn9b { background-color: rgb(66, 133, 244); }

.misTTe { transform: translate(0px, 0px); }

@media screen and (min-width: 481px) {
  .Mh0NNb { min-width: 288px; max-width: 568px; border-radius: 2px; }
  .Mp2Z0b { left: 24px; margin-right: 24px; right: auto; }
  .VcC8Fc { left: 50%; right: auto; transform: translate(-50%, 100%); }
  .Mp2Z0b.misTTe { bottom: 24px; }
  .VcC8Fc.misTTe { bottom: 0px; transform: translate(-50%, 0px); }
  .M6tHv { padding: 0px; }
  .aGJE1b { padding-right: 24px; }
}

@media screen and (max-width: 480px) {
  .xbgI6e .aGJE1b, .xbgI6e .x95qze { padding-bottom: 24px; padding-top: 24px; }
}

@media screen and (min-width: 481px) and (max-width: 568px) {
  .Mh0NNb { max-width: 90%; }
}

@media screen and (min-width: 569px) {
  .Mh0NNb { max-width: 568px; }
}

.XzbSje { border: 1px solid transparent; border-radius: var(--dt-corner-banner,.25rem); box-sizing: border-box; background: var(--dt-background,#fff); color: var(--dt-on-background,rgb(60,64,67)); display: flex; padding: 0.6875rem 0.4375rem 0.6875rem 0.9375rem; transition: height 0.25s cubic-bezier(0, 0, 0.2, 1) 0s, margin 0.25s cubic-bezier(0, 0, 0.2, 1) 0s; user-select: text; }

.vhoiae .XzbSje, .X9XeLb .XzbSje, .cWKK1c .XzbSje, .aJfoSc .XzbSje, .TOb6Ze .XzbSje { padding-bottom: 0.8125rem; padding-top: 0.8125rem; }

.XzbSje.fs1v2 { padding-right: 0.9375rem; }

.XzbSje:not(.eO2Zfd) { border-width: 0px; height: 0px; margin: 0px; min-height: 0px; padding: 0px; transition: height 0.25s cubic-bezier(0, 0, 0.2, 1) 0s, margin 0.25s cubic-bezier(0, 0, 0.2, 1) 0s, visibility 0.25s step-end 0s; visibility: hidden; }

.XzbSje.hECuDf { border-radius: 0px; }

.XzbSje.UkbGab { padding: 0.4375rem 0.4375rem 0.4375rem 0.9375rem; }

.mLhC9c { height: 0px; opacity: 0; position: fixed; top: -5000px; width: 0px; }

.EPX8Dc { box-sizing: border-box; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; margin-right: 1rem; max-height: 8rem; max-width: 8rem; }

.EPX8Dc.bkJe8c { -webkit-box-align: center; align-items: center; fill: currentcolor; height: 1.25rem; width: 1.25rem; }

.EPX8Dc.hECuDf { margin-left: 0.5rem; margin-right: 1.5rem; }

.EPX8Dc.MELUue { margin: 0.5rem 1rem 0.5rem 0.5rem; }

.R7nqif { fill: currentcolor; font-weight: 500; margin-left: 0.25em; }

.eZZewe.vKmmhc { -webkit-box-align: center; align-items: center; display: flex; height: 2.25rem; -webkit-box-pack: center; justify-content: center; margin: 0px; padding: 0px; width: 2.25rem; }

.eZZewe.vKmmhc.UkbGab { height: 1.75rem; width: 1.75rem; }

.SPs1Af { display: flex; }

.SPs1Af.vKmmhc.UkbGab { height: 1.125rem; width: 1.125rem; }

.zRDX4b { z-index: 6000; }

.le1PVb { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); align-self: center; -webkit-box-flex: 1; flex: 1 1 auto; margin-bottom: 0.75rem; }

.le1PVb:not(.fs1v2) { margin-right: 0.5rem; }

.xUlw3b { font: var(--dt-headline-6-font,400 1.125rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-headline-6-spacing,0); flex-basis: 100%; margin-bottom: 0.25rem; }

.DGjo0e { font-style: ; font-variant-ligatures: ; font-variant-caps: ; font-variant-numeric: ; font-variant-east-asian: ; font-variant-alternates: ; font-stretch: ; font-size: ; line-height: ; font-family: ; font-optical-sizing: ; font-kerning: ; font-feature-settings: ; font-variation-settings: ; letter-spacing: var(--dt-title-small-spacing,.0178571429em); display: inline-flex; -webkit-box-flex: 0; flex: 0 1 auto; font-weight: 500; padding-right: 0.5ch; }

.nuPcl { -webkit-box-align: center; align-items: center; align-self: flex-end; animation: 0.2s linear 0s 1 normal backwards running driveBannerActionsEntrance; box-sizing: border-box; display: flex; -webkit-box-flex: 1; flex: 1 0 auto; height: 1.25rem; -webkit-box-pack: end; justify-content: flex-end; margin-bottom: 0.75rem; }

@-webkit-keyframes driveBannerActionsEntrance { 
  0% { opacity: 0; visibility: hidden; }
}

@keyframes driveBannerActionsEntrance { 
  0% { opacity: 0; visibility: hidden; }
}

.vhoiae .nuPcl, .X9XeLb .nuPcl, .cWKK1c .nuPcl, .aJfoSc .nuPcl, .TOb6Ze .nuPcl, .nuPcl.UkbGab { height: 1.25rem; }

.nuPcl.WGEhue { width: 100%; }

.kYqbf { margin-left: 0.25rem; }

.kYqbf.vKmmhc.UkbGab { height: 1.75rem; }

.XzbSje.cEsmJb .nuPcl { -webkit-box-flex: 0; flex: 0 0 auto; }

.iLpyV { -webkit-box-align: center; align-items: center; box-sizing: border-box; display: flex; -webkit-box-flex: 0; flex: 0 0 auto; height: 1.25rem; padding: 0.125rem; }

.vhoiae .iLpyV, .X9XeLb .iLpyV, .cWKK1c .iLpyV, .aJfoSc .iLpyV, .TOb6Ze .iLpyV, .XzbSje.UkbGab .iLpyV { height: 1.25rem; }

.br9Wvc { box-sizing: border-box; -webkit-box-flex: 1; flex: 1 1 auto; flex-wrap: wrap; max-width: 100%; }

.Dsuz9e { align-self: center; align-content: space-between; display: flex; -webkit-box-flex: 1; flex: 1 1 100%; flex-wrap: wrap; margin-bottom: -0.75rem; min-height: 2rem; }

.vhoiae .Dsuz9e, .X9XeLb .Dsuz9e, .cWKK1c .Dsuz9e, .aJfoSc .Dsuz9e, .TOb6Ze .Dsuz9e, .Dsuz9e.UkbGab { min-height: 2rem; }

.Dsuz9e.MELUue { padding: 0.5rem 0.5rem 0.75rem; }

.Dsuz9e.MELUue.wg2eAc { padding-bottom: 0.25rem; }

.Dsuz9e.WGEhue { align-self: stretch; }

.vbK9Ff { display: flex; -webkit-box-flex: 1; flex: 1 1 100%; }

.XzbSje.eO2Zfd .nuPcl, .XzbSje.eO2Zfd .br9Wvc, .XzbSje.eO2Zfd .EPX8Dc { transition: opacity 50ms linear 0.2s; }

.XzbSje:not(.eO2Zfd) .nuPcl, .XzbSje:not(.eO2Zfd) .br9Wvc, .XzbSje:not(.eO2Zfd) .EPX8Dc { opacity: 0; transition: opacity 50ms linear 0s; }

.XzbSje.T3YfFf, .XzbSje.T3YfFf .nuPcl, .XzbSje.T3YfFf .br9Wvc, .XzbSje.T3YfFf .EPX8Dc { transition-duration: 1ms; }

.XzbSje.w8ecmf.VLrnY { background: var(--dt-neutral-container,rgb(241,243,244)); border-color: var(--dt-neutral-container,rgb(241,243,244)); color: var(--dt-on-neutral-container,rgb(60,64,67)); }

.XzbSje.w8ecmf.I5JVbf { border-color: var(--dt-neutral-outline,rgb(60,64,67)); color: var(--dt-on-neutral-container,rgb(60,64,67)); }

.XzbSje.w8ecmf.eJxL0c { background: var(--dt-neutral,rgb(60,64,67)); border-color: var(--dt-neutral,rgb(60,64,67)); color: var(--dt-on-neutral,#fff); }

.XzbSje.AVUQbb.VLrnY { background: var(--dt-primary-container,rgb(232,240,254)); border-color: var(--dt-primary-container,rgb(232,240,254)); color: var(--dt-on-primary-container,rgb(60,64,67)); }

.XzbSje.AVUQbb.I5JVbf { border-color: var(--dt-primary-outline,rgb(24,90,188)); color: var(--dt-on-primary-container,rgb(60,64,67)); }

.XzbSje.AVUQbb.eJxL0c { background: var(--dt-primary,rgb(26,115,232)); border-color: var(--dt-primary,rgb(26,115,232)); color: var(--dt-on-primary,#fff); }

.XzbSje.S9cmWe.VLrnY { background: var(--dt-warning-container,rgb(254,247,224)); border-color: var(--dt-warning-container,rgb(254,247,224)); color: var(--dt-on-warning-container,rgb(60,64,67)); }

.XzbSje.S9cmWe.I5JVbf { border-color: var(--dt-warning-outline,rgb(234,134,0)); color: var(--dt-on-warning-container,rgb(60,64,67)); }

.XzbSje.S9cmWe.eJxL0c { background: var(--dt-warning,rgb(249,171,0)); border-color: var(--dt-warning,rgb(249,171,0)); color: var(--dt-on-warning,rgb(32,33,36)); }

.XzbSje.m586Kb.VLrnY { background: var(--dt-error-container,rgb(252,232,230)); border-color: var(--dt-error-container,rgb(252,232,230)); color: var(--dt-on-error-container,rgb(60,64,67)); }

.XzbSje.m586Kb.I5JVbf { border-color: var(--dt-error-outline,rgb(179,20,18)); color: var(--dt-on-error-container,rgb(60,64,67)); }

.XzbSje.m586Kb.eJxL0c { background: var(--dt-error,rgb(217,48,37)); border-color: var(--dt-error,rgb(217,48,37)); color: var(--dt-on-error,#fff); }

.XzbSje.aUai5e.VLrnY { background: var(--dt-tertiary-container,rgb(230,244,234)); border-color: var(--dt-tertiary-container,rgb(230,244,234)); color: var(--dt-on-tertiary-container,rgb(60,64,67)); }

.XzbSje.aUai5e.I5JVbf { border-color: var(--dt-tertiary-outline,rgb(19,115,51)); color: var(--dt-on-tertiary-container,rgb(60,64,67)); }

.XzbSje.aUai5e.eJxL0c { background: var(--dt-tertiary,rgb(24,128,56)); border-color: var(--dt-tertiary,rgb(24,128,56)); color: var(--dt-on-tertiary,#fff); }

.R7nqif.w8ecmf.VLrnY, .R7nqif.w8ecmf.I5JVbf { color: var(--dt-neutral-container-link,rgb(25,103,210)); }

.R7nqif.w8ecmf.eJxL0c { color: var(--dt-neutral-link,#fff); }

.R7nqif.AVUQbb.VLrnY, .R7nqif.AVUQbb.I5JVbf { color: var(--dt-primary-container-link,rgb(25,103,210)); }

.R7nqif.AVUQbb.eJxL0c { color: var(--dt-primary-link,#fff); }

.R7nqif.S9cmWe.VLrnY, .R7nqif.S9cmWe.I5JVbf { color: var(--dt-warning-container-link,rgb(60,64,67)); }

.R7nqif.S9cmWe.eJxL0c { color: var(--dt-warning-link,rgb(60,64,67)); }

.R7nqif.m586Kb.VLrnY, .R7nqif.m586Kb.I5JVbf { color: var(--dt-error-container-link,rgb(197,34,31)); }

.R7nqif.m586Kb.eJxL0c { color: var(--dt-error-link,#fff); }

.R7nqif.aUai5e.VLrnY, .R7nqif.aUai5e.I5JVbf { color: var(--dt-tertiary-container-link,rgb(19,115,51)); }

.R7nqif.aUai5e.eJxL0c { color: var(--dt-tertiary-link,#fff); }

.EPX8Dc.w8ecmf.VLrnY, .EPX8Dc.w8ecmf.I5JVbf { color: var(--dt-neutral-container-icon,rgb(60,64,67)); }

.EPX8Dc.w8ecmf.eJxL0c { color: var(--dt-neutral-icon,#fff); }

.EPX8Dc.AVUQbb.VLrnY, .EPX8Dc.AVUQbb.I5JVbf { color: var(--dt-primary-container-icon,rgb(25,103,210)); }

.EPX8Dc.AVUQbb.eJxL0c { color: var(--dt-primary-icon,#fff); }

.EPX8Dc.S9cmWe.VLrnY, .EPX8Dc.S9cmWe.I5JVbf { color: var(--dt-warning-container-icon,rgb(60,64,67)); }

.EPX8Dc.S9cmWe.eJxL0c { color: var(--dt-warning-icon,rgb(60,64,67)); }

.EPX8Dc.m586Kb.VLrnY, .EPX8Dc.m586Kb.I5JVbf { color: var(--dt-error-container-icon,rgb(197,34,31)); }

.EPX8Dc.m586Kb.eJxL0c { color: var(--dt-error-icon,#fff); }

.EPX8Dc.aUai5e.VLrnY, .EPX8Dc.aUai5e.I5JVbf { color: var(--dt-tertiary-container-icon,rgb(19,115,51)); }

.EPX8Dc.aUai5e.eJxL0c { color: var(--dt-tertiary-icon,#fff); }

.vhoiae .grsXwb, .X9XeLb .grsXwb, .cWKK1c .grsXwb, .aJfoSc .grsXwb, .TOb6Ze .grsXwb { width: 20px; height: 20px; }

.llhEMd { transition: opacity 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0.15s; background-color: rgba(0, 0, 0, 0.5); inset: 0px; opacity: 0; position: fixed; z-index: 5000; }

.llhEMd.iWO5td { transition: opacity 0.05s cubic-bezier(0.4, 0, 0.2, 1) 0s; opacity: 1; }

.mjANdc { transition: transform 0.4s cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 0.4s cubic-bezier(0.4, 0, 0.2, 1) 0s; -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: vertical; flex-direction: column; inset: 0px; padding: 0px 5%; position: absolute; }

.x3wWge, .ONJhl { display: block; height: 3em; }

.eEPege > .x3wWge, .eEPege > .ONJhl { -webkit-box-flex: 1; flex-grow: 1; }

.J9Nfi { flex-shrink: 1; max-height: 100%; }

.g3VIld { -webkit-box-align: stretch; align-items: stretch; display: flex; -webkit-box-orient: vertical; flex-direction: column; transition: transform 0.225s cubic-bezier(0, 0, 0.2, 1) 0s, -webkit-transform 0.225s cubic-bezier(0, 0, 0.2, 1) 0s; position: relative; background-color: rgb(255, 255, 255); border-radius: 2px; box-shadow: rgba(0, 0, 0, 0.24) 0px 12px 15px 0px; max-width: 24em; outline: transparent solid 1px; overflow: hidden; }

.vcug3d .g3VIld { padding: 0px; }

.g3VIld.kdCdqc { transition: transform 0.15s cubic-bezier(0.4, 0, 1, 1) 0s, -webkit-transform 0.15s cubic-bezier(0.4, 0, 1, 1) 0s; }

.Up8vH.CAwICe { transform: scale(0.8); }

.Up8vH.kdCdqc { transform: scale(0.9); }

.E4P6x.CAwICe, .E4P6x.kdCdqc { transform: translateY(50%); }

.vDc8Ic.CAwICe { transform: scale(0.8) translateY(100%); }

.XIJ9Ac > .x3wWge, .XIJ9Ac > .ONJhl, .HhoEBe > .x3wWge { -webkit-box-flex: 1; flex-grow: 1; }

.HhoEBe > .ONJhl { -webkit-box-flex: 2; flex-grow: 2; }

.Nevtdc > .x3wWge { -webkit-box-flex: 0; flex-grow: 0; }

.Nevtdc > .ONJhl, .t8Vtv > .x3wWge { -webkit-box-flex: 1; flex-grow: 1; }

.t8Vtv > .g3VIld { -webkit-box-flex: 2; flex-grow: 2; }

.t8Vtv > .ONJhl { -webkit-box-flex: 1; flex-grow: 1; }

.vcug3d { -webkit-box-align: stretch; align-items: stretch; padding: 0px; }

.vcug3d > .g3VIld { -webkit-box-flex: 2; flex-grow: 2; border-radius: 0px; left: 0px; right: 0px; max-width: 100%; }

.vcug3d > .ONJhl, .vcug3d > .x3wWge { -webkit-box-flex: 0; flex-grow: 0; height: 0px; }

.tOrNgd { display: flex; flex-shrink: 0; font: 500 20px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 24px 24px 20px; }

.vcug3d .tOrNgd { display: none; }

.TNczib { -webkit-box-pack: justify; justify-content: space-between; flex-shrink: 0; box-shadow: rgba(0, 0, 0, 0.24) 0px 3px 4px 0px; background-color: rgb(69, 90, 100); color: white; display: none; font: 500 20px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.vcug3d .TNczib { display: flex; }

.PNenzf { -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; overflow: hidden; overflow-wrap: break-word; }

.TNczib .PNenzf { margin: 16px 0px; }

.VY7JQd { height: 0px; }

.TNczib .VY7JQd, .tOrNgd .bZWIgd { display: none; }

.R6Lfte .Wtw8H { flex-shrink: 0; display: block; margin: -12px -6px 0px 0px; }

.PbnGhe { -webkit-box-flex: 2; flex-grow: 2; flex-shrink: 2; display: block; font: 400 14px / 20px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 0px 24px; overflow-y: auto; }

.Whe8ub .PbnGhe { padding-top: 24px; }

.hFEqNb .PbnGhe { padding-bottom: 24px; }

.vcug3d .PbnGhe { padding: 16px; }

.XfpsVe { display: flex; flex-shrink: 0; -webkit-box-pack: end; justify-content: flex-end; padding: 24px 24px 16px; }

.vcug3d .XfpsVe { display: none; }

.OllbWe { -webkit-box-pack: end; justify-content: flex-end; display: none; }

.vcug3d .OllbWe { display: flex; -webkit-box-align: start; align-items: flex-start; margin: 0px 16px; }

.kHssdc.O0WRkf.C0oVfc, .XfpsVe .O0WRkf.C0oVfc { min-width: 64px; }

.kHssdc + .kHssdc { margin-left: 8px; }

.TNczib .kHssdc { color: rgb(255, 255, 255); margin-top: 10px; }

.TNczib .Wtw8H { margin: 4px 24px 4px 0px; }

.TNczib .kHssdc.u3bW4e, .TNczib .Wtw8H.u3bW4e { background-color: rgba(204, 204, 204, 0.25); }

.TNczib .kHssdc > .Vwe4Vb, .TNczib .Wtw8H > .VTBa7b { background-image: radial-gradient(circle farthest-side, rgba(255, 255, 255, 0.3), rgba(255, 255, 255, 0.3) 80%, rgba(255, 255, 255, 0) 100%); }

.TNczib .kHssdc.RDPZE, .TNczib .Wtw8H.RDPZE { color: rgba(255, 255, 255, 0.5); fill: rgba(255, 255, 255, 0.5); }

.VUI3Tc { overflow: auto; }

.nkvGQ { display: none; }

.nkvGQ.O9rvMd { display: block; position: absolute; top: 0px; background-color: black; opacity: 0.4; height: 100%; width: 100%; z-index: 2000; }

.wrPvic { border-radius: 8px; height: auto; max-width: 640px; min-height: 570px; overflow: visible; width: 640px; }

.wrPvic .qRUolc { padding-bottom: 15px; padding-top: 20px; }

.wrPvic .J9fJmf { -webkit-box-align: center; align-items: center; padding-bottom: 20px; }

.wrPvic .oJeWuf { overflow-y: visible; }

.XKAX7, .dEW8tb { padding: 0px 16px; text-transform: none; font: var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-medium-spacing,.00625em); }

.XKAX7 { color: var(--dt-primary,rgb(26,115,232)); margin-right: 16px; min-width: 50px; }

.XKAX7:hover { background-color: var(--dt-primary-container,rgb(232,240,254)); }

.dEW8tb { background-color: var(--dt-primary,rgb(26,115,232)); border-radius: 4px; box-shadow: none; }

.dEW8tb[disabled] { background-color: rgba(153, 153, 153, 0.1); }

.dEW8tb:not([disabled]):hover { background-color: var(--dt-primary-action-state-layer,rgb(25,103,210)); border-radius: 4px; box-shadow: 0px 1px 2px 0px; }

.XKAX7 .snByac, .dEW8tb .snByac { margin: 8px 16px; }

.Xs9kmd { -webkit-box-flex: 1; flex-grow: 1; margin-left: 2px; }

.oqO1sd { color: var(--dt-on-surface-variant,rgb(95,99,104)); margin-bottom: 16px; margin-top: 8px; font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); }

.fE2C5b { -webkit-box-align: center; align-items: center; display: flex; }

.fE2C5b .ZaiL8e { fill: var(--dt-primary,rgb(26,115,232)); height: 24px; padding-right: 16px; width: 24px; }

.BrvSpf { font: var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-title-large-spacing,0); color: var(--dt-on-surface,rgb(60,64,67)); }

.b8odnb { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; height: 100%; position: relative; width: 100%; }

.zzuIoc, .XEMjs { width: 100%; }

.OxFvPe { border: 1px solid var(--dt-outline,rgb(128,134,139)); border-radius: 100px; display: inline-block; font-size: 14px; height: 32px; max-width: 550px; padding-left: 15px; padding-right: 15px; }

.ZpZNmb { -webkit-box-align: center; align-items: center; display: flex; height: 100%; }

.MuyDde { overflow-x: hidden; padding-left: 10px; text-overflow: ellipsis; }

.URwq { color: var(--dt-error,rgb(217,48,37)); display: none; -webkit-box-flex: 1; flex-grow: 1; flex-shrink: 1; margin-bottom: 16px; margin-top: 8px; font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); }

.URwq.McD6Rc { display: block; }

.qzWk0c { -webkit-box-align: center; align-items: center; background-color: var(--dt-primary-container,rgb(232,240,254)); border-radius: 8px; display: flex; margin-top: 8px; }

.MeX0je { color: var(--dt-on-primary-container,rgb(60,64,67)); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); }

.b8odnb.uNaCce .qzWk0c { background-color: var(--dt-tertiary-container,rgb(230,244,234)); }

.b8odnb.uNaCce .MeX0je { display: none; }

.v7tbof { display: none; color: var(--dt-tertiary,rgb(24,128,56)); font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); }

.b8odnb.uNaCce .v7tbof { display: block; }

.CzZ0kd { margin: 16px 0px 12px; }

.D1rc6d { border-radius: 8px; left: 2px; position: absolute; right: unset; top: 0px; }

.TP8uyc { box-sizing: border-box; color: var(--dt-background,#fff); transition: background 0.25s linear 0s, color 0.25s linear 0s; }

.TP8uyc.aQE9pc { background: rgb(248, 249, 250); position: relative; }

.TP8uyc.aQE9pc::after { border-radius: 100px; border: 2px solid transparent; box-sizing: border-box; content: ""; display: block; height: 100%; left: 0px; pointer-events: none; position: absolute; top: 0px; width: 100%; }

.AsSTTb { -webkit-box-align: center; place-items: center; background: rgb(239, 239, 239); border-radius: 100px; box-sizing: border-box; display: flex; font-family: "Google Sans"; font-size: 1rem; -webkit-box-pack: center; justify-content: center; position: relative; text-align: center; text-transform: uppercase; -webkit-box-flex: 0; flex: 0 0 auto; text-overflow: ellipsis; white-space: nowrap; }

.AsSTTb.EwXqJf { height: 2.75rem; width: 2.75rem; }

.AsSTTb.NWlIHc { height: 2.5rem; width: 2.5rem; }

.AsSTTb.nsKVp { font-size: 1.125rem; height: 2.25rem; width: 2.25rem; }

.AsSTTb.GND07b { font-size: 1rem; height: 2rem; width: 2rem; }

.AsSTTb.SjheHf { font-size: 1rem; height: 1.5rem; width: 1.5rem; }

.AsSTTb.HHWuM { font-size: 0.75rem; height: 1.25rem; width: 1.25rem; }

.AsSTTb.Ppq72 { font-size: 0.75rem; height: 1rem; width: 1rem; }

.AsSTTb.aQE9pc { background: rgb(248, 249, 250); }

.lezq { border-radius: inherit; box-sizing: border-box; letter-spacing: -0.035ch; margin-top: 0.035ex; opacity: 0.75; }

.lezq.EwXqJf { font-size: 1.75rem; }

.lezq.NWlIHc { font-size: 1.5rem; }

.lezq.nsKVp { font-size: 1.25rem; }

.lezq.GND07b { font-size: 1.125rem; }

.lezq.SjheHf { font-size: 1rem; }

.HYmxfb { -webkit-box-align: center; align-items: center; border: 1px solid transparent; border-radius: inherit; box-sizing: border-box; display: inline-flex; height: 100%; -webkit-box-pack: center; justify-content: center; width: 100%; }

.HYmxfb.TVtO8d { background: var(--dt-primary,rgb(26,115,232)); }

.HYmxfb.SGdsQe { background: rgb(30, 142, 62); }

.HYmxfb.uUAVm { background: rgb(242, 153, 0); }

.HYmxfb.X7pJl { background: rgb(232, 113, 10); }

.HYmxfb.RnwtS { background: var(--dt-error,rgb(217,48,37)); }

.HYmxfb.nhV17d { background: rgb(229, 37, 146); }

.HYmxfb.usAlUd { background: rgb(147, 52, 230); }

.HYmxfb.kuBvP { background: rgb(18, 181, 203); }

.HYmxfb.TLMa7e { color: var(--dt-background,#fff); background: rgb(189, 193, 198); }

.GOZObd { background: var(--dt-background,#fff); border-radius: inherit; box-sizing: border-box; color: var(--dt-outline-variant,rgb(218,220,224)); height: 100%; transition: color 0.25s linear 0s; width: 100%; }

.SdHJPc { border-radius: inherit; box-sizing: border-box; height: 100%; width: 100%; }

.uS40rb { border-radius: inherit; box-sizing: border-box; height: inherit; width: inherit; }

.uS40rb.pyzYhb { height: 1rem; width: 1rem; }

.uS40rb.pyzYhb.EwXqJf { height: 1.75rem; width: 1.75rem; }

.uS40rb.pyzYhb.NWlIHc { height: 1.5rem; width: 1.5rem; }

.uS40rb.pyzYhb.nsKVp { height: 1.25rem; width: 1.25rem; }

.uS40rb.pyzYhb.GND07b { height: 1.125rem; width: 1.125rem; }

.bhxwjd { align-items: center; background-color: transparent; display: flex; -webkit-box-flex: 1; flex-grow: 1; max-width: 100%; min-height: 37px; }

.YMNIz { overflow: hidden; width: 100%; }

.YMNIz::before { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; color: var(--dt-on-surface-variant,#5f6368); content: attr(data-before-input); outline: transparent solid 1px; white-space: pre-wrap; word-break: break-all; }

.YMNIz::after { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; color: var(--dt-on-surface-variant,#5f6368); content: attr(data-after-input); outline: transparent solid 1px; white-space: pre-wrap; word-break: break-all; }

.zeumMd { letter-spacing: 0.0142857em; font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; font-weight: 400; line-height: 1.25rem; background-color: transparent; border: none; caret-color: var(--dt-primary,#1a73e8); color: var(--dt-on-surface,#3c4043); width: 1px; min-height: 1em; outline: transparent solid 1px; overflow: auto; padding: 0px; white-space: nowrap; }

.zeumMd.d2j1H { margin-right: -100%; padding-right: 100%; }

.zeumMd::-webkit-scrollbar { display: none; }

.zeumMd.NDUvFb { height: 0px; position: absolute; white-space: pre; visibility: hidden; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-qrOfGf { position: absolute; top: 50%; height: 48px; left: 50%; width: 48px; transform: translate(-50%, -50%); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { border: none; display: inline-flex; position: relative; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; box-sizing: border-box; padding: 0px; outline: none; cursor: pointer; appearance: none; background: none; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-f2wwtd { height: 18px; width: 18px; font-size: 18px; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-qrOfGf { width: 26px; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-f2wwtd { fill: currentcolor; color: inherit; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { top: 0px; left: 0px; width: 100%; height: 100%; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000)); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob { position: absolute; box-sizing: content-box; width: 100%; height: 100%; overflow: hidden; }

.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgba(0, 0, 0, 0.54); }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: rgb(0, 0, 0); }

.VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgba(0, 0, 0, 0.54); }

.VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgba(0, 0, 0, 0.62); }

.VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgba(0, 0, 0, 0.87); }

.VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { width: 20px; height: 20px; font-size: 20px; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-f2wwtd { height: 18px; width: 18px; font-size: 18px; }

.VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-UbuQg { width: 18px; height: 18px; font-size: 18px; }

.VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { margin-left: 4px; margin-right: -4px; }

[dir="rtl"] .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc[dir="rtl"] { margin-left: -4px; margin-right: 4px; }

.VfPpkd-Zr1Nwf-OWXEXe-UbuQg { margin-left: 4px; margin-right: -4px; }

[dir="rtl"] .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .VfPpkd-Zr1Nwf-OWXEXe-UbuQg[dir="rtl"] { margin-left: -4px; margin-right: 4px; }

.VfPpkd-XPtOyb { border-radius: 16px; background-color: rgb(224, 224, 224); color: rgba(0, 0, 0, 0.87); -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-body2-font-size,.875rem); line-height: var(--mdc-typography-body2-line-height,1.25rem); font-weight: var(--mdc-typography-body2-font-weight,400); letter-spacing: var(--mdc-typography-body2-letter-spacing,.0178571429em); text-decoration: var(--mdc-typography-body2-text-decoration,inherit); text-transform: var(--mdc-typography-body2-text-transform,inherit); height: 32px; position: relative; display: inline-flex; -webkit-box-align: center; align-items: center; box-sizing: border-box; padding: 0px 12px; border-width: 0px; outline: none; cursor: pointer; appearance: none; }

.VfPpkd-XPtOyb .VfPpkd-v1cqY { border-radius: 16px; }

.VfPpkd-XPtOyb:hover { color: rgba(0, 0, 0, 0.87); }

.VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, .VfPpkd-XPtOyb .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { margin-left: -4px; margin-right: 4px; }

[dir="rtl"] .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, [dir="rtl"] .VfPpkd-XPtOyb .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce), .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir="rtl"], .VfPpkd-XPtOyb .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir="rtl"] { margin-left: 4px; margin-right: -4px; }

.VfPpkd-XPtOyb .VfPpkd-BFbNVe-bF1uUb { width: 100%; height: 100%; top: 0px; left: 0px; }

.VfPpkd-XPtOyb:hover { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-XPtOyb .VfPpkd-lrT0x { position: absolute; top: 50%; height: 48px; left: 0px; right: 0px; transform: translateY(-50%); }

.VfPpkd-XPtOyb-OWXEXe-SNIJTd { transition: opacity 75ms cubic-bezier(0.4, 0, 0.2, 1) 0s, width 0.15s cubic-bezier(0, 0, 0.2, 1) 0s, padding 0.1s linear 0s, margin 0.1s linear 0s; opacity: 0; }

.VfPpkd-WX5mde { text-overflow: ellipsis; overflow: hidden; }

.VfPpkd-TfeOUb { white-space: nowrap; }

.VfPpkd-Zr1Nwf { border-radius: 50%; outline: none; vertical-align: middle; }

.VfPpkd-PvL5qd { height: 20px; }

.VfPpkd-PvL5qd-Jt5cK { transition: stroke-dashoffset 0.15s cubic-bezier(0.4, 0, 0.6, 1) 50ms; stroke-width: 2px; stroke-dashoffset: 29.7833; stroke-dasharray: 29.7833; }

.VfPpkd-rXoKne-JIbuQc:focus { outline: none; }

.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd-Jt5cK { stroke-dashoffset: 0; }

.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { position: relative; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgba(98, 0, 238, 0.54); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb .VfPpkd-PvL5qd-Jt5cK { stroke: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb-OWXEXe-gk6SMd { background-color: var(--mdc-theme-surface,#fff); }

.VfPpkd-PvL5qd-OAU7Vd { width: 0px; height: 20px; transition: width 0.15s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd-OAU7Vd { width: 20px; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { transition: opacity 75ms linear -50ms; opacity: 1; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc + .VfPpkd-PvL5qd { transition: opacity 75ms linear 80ms; opacity: 0; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc + .VfPpkd-PvL5qd .VfPpkd-PvL5qd-OAU7Vd { transition: width 0ms ease 0s; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { opacity: 0; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc + .VfPpkd-PvL5qd { width: 0px; opacity: 1; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { width: 0px; opacity: 0; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-yOOK0 .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc + .VfPpkd-PvL5qd { width: 20px; }

.VfPpkd-XPtOyb { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-XPtOyb .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb .VfPpkd-v1cqY::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-XPtOyb .VfPpkd-v1cqY::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-XPtOyb .VfPpkd-v1cqY::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d .VfPpkd-v1cqY::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d .VfPpkd-v1cqY::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-v1cqY::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-v1cqY::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-v1cqY::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-XPtOyb .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb .VfPpkd-v1cqY::after { top: -50%; left: -50%; width: 200%; height: 200%; }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d .VfPpkd-v1cqY::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-XPtOyb .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb .VfPpkd-v1cqY::after { background-color: var(--mdc-ripple-color,rgba(0,0,0,.87)); }

.VfPpkd-XPtOyb:hover .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb:focus-within .VfPpkd-v1cqY::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-XPtOyb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-XPtOyb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-XPtOyb.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-XPtOyb .VfPpkd-v1cqY { position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; pointer-events: none; overflow: hidden; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-selected-opacity,.08); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-hover-opacity,.12); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before, .VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus-within .VfPpkd-v1cqY::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.2); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.2); }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-X7AZM .VfPpkd-XPtOyb.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.2); }

@-webkit-keyframes mdc-chip-entry { 
  0% { transform: scale(0.8); opacity: 0.4; }
  100% { transform: scale(1); opacity: 1; }
}

@keyframes mdc-chip-entry { 
  0% { transform: scale(0.8); opacity: 0.4; }
  100% { transform: scale(1); opacity: 1; }
}

.VfPpkd-XPtOyb-FCjw3e { padding: 4px; display: flex; flex-wrap: wrap; box-sizing: border-box; }

.VfPpkd-XPtOyb-FCjw3e .VfPpkd-XPtOyb { margin: 4px; }

.VfPpkd-XPtOyb-FCjw3e .VfPpkd-XPtOyb-OWXEXe-dgl2Hf { margin-top: 8px; margin-bottom: 8px; }

.VfPpkd-XPtOyb-FCjw3e-OWXEXe-YPqjbf .VfPpkd-XPtOyb { animation: 0.1s cubic-bezier(0, 0, 0.2, 1) 0s 1 normal none running mdc-chip-entry; }

.P2wJPb { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; z-index: 0; color: var(--gm-chip-ink-color,rgb(95,99,104)); }

.P2wJPb.VfPpkd-XPtOyb-OWXEXe-SNIJTd { transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s, opacity 75ms cubic-bezier(0.4, 0, 0.2, 1) 0s, width 0.15s cubic-bezier(0, 0, 0.2, 1) 0s, padding 0.1s linear 0s, margin 0.1s linear 0s; }

.P2wJPb .VfPpkd-v1cqY::before, .P2wJPb .VfPpkd-v1cqY::after { z-index: -1; }

.P2wJPb .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(95, 99, 104); }

.P2wJPb .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color,rgb(95,99,104)); }

.P2wJPb .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(95, 99, 104); }

.P2wJPb .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(95, 99, 104); }

.P2wJPb .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(95, 99, 104); }

.P2wJPb .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color,rgb(95,99,104)); }

.P2wJPb:hover, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus, .P2wJPb:active { color: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.P2wJPb:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(32, 33, 36); }

.P2wJPb:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.P2wJPb:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(32, 33, 36); }

.P2wJPb:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(32, 33, 36); }

.P2wJPb:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(32, 33, 36); }

.P2wJPb:hover .VfPpkd-PvL5qd-Jt5cK, .P2wJPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK, .P2wJPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK, .P2wJPb:active .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd { background-color: var(--gm-chip-container-color,rgb(232,240,254)); color: var(--gm-chip-ink-color,rgb(25,103,210)); border-color: var(--gm-chip-outline-color--stateful,rgb(23,78,166)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(25, 103, 210); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color,rgb(25,103,210)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(25, 103, 210); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(25, 103, 210); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(25, 103, 210); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color,rgb(25,103,210)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active { color: var(--gm-chip-ink-color--stateful,rgb(23,78,166)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(23, 78, 166); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color--stateful,rgb(23,78,166)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(23, 78, 166); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(23, 78, 166); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(23, 78, 166); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-PvL5qd-Jt5cK, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color--stateful,rgb(23,78,166)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::before, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::after { background-color: var(--gm-chip-state-color,rgb(25,103,210)); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-v1cqY::before, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before, .P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after { transition: opacity 0.15s linear 0s; }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.P2wJPb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.YfmZeb { background-color: var(--gm-chip-container-color,transparent); border-style: solid; padding-right: 15px; padding-left: 15px; border-width: 1px; border-color: var(--gm-chip-outline-color,rgb(218,220,224)); }

.YfmZeb .VfPpkd-v1cqY { top: -1px; left: -1px; border: 1px solid transparent; }

.YfmZeb .VfPpkd-v1cqY::before, .YfmZeb .VfPpkd-v1cqY::after { background-color: var(--gm-chip-state-color,rgb(60,64,67)); }

.YfmZeb:hover .VfPpkd-v1cqY::before, .YfmZeb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.YfmZeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before, .YfmZeb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.YfmZeb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after { transition: opacity 0.15s linear 0s; }

.YfmZeb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.YfmZeb.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.YfmZeb:focus, .YfmZeb.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe { border-color: var(--gm-chip-outline-color--stateful,rgb(32,33,36)); }

.YfmZeb:active { box-shadow: none; }

.YfmZeb:active .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd { padding-right: 16px; padding-left: 16px; border-width: 0px; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY { top: 0px; left: 0px; border: 0px solid transparent; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover { box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus, .YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe { padding-right: 15px; padding-left: 15px; border-width: 1px; }

.YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus .VfPpkd-v1cqY, .YfmZeb.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe .VfPpkd-v1cqY { top: -1px; left: -1px; border: 1px solid transparent; }

.MUK9yc { background-color: var(--gm-chip-container-color,#fff); padding-right: 16px; padding-left: 16px; border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.MUK9yc .VfPpkd-v1cqY::before, .MUK9yc .VfPpkd-v1cqY::after { background-color: var(--gm-chip-state-color,rgb(60,64,67)); }

.MUK9yc:hover .VfPpkd-v1cqY::before, .MUK9yc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.MUK9yc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before, .MUK9yc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.MUK9yc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after { transition: opacity 0.15s linear 0s; }

.MUK9yc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.MUK9yc.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.MUK9yc .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.MUK9yc:hover { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.MUK9yc:hover .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.MUK9yc:active { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; }

.MUK9yc:active .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.tTvXye { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; padding-right: 11px; padding-left: 11px; border-width: 1px; }

.tTvXye .VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { width: 20px; height: 20px; font-size: 20px; }

.tTvXye.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, .tTvXye .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { margin-left: -3px; margin-right: 8px; }

[dir="rtl"] .tTvXye.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, [dir="rtl"] .tTvXye .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce), .tTvXye.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir="rtl"], .tTvXye .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir="rtl"] { margin-left: 8px; margin-right: -3px; }

.tTvXye .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { margin-left: 8px; margin-right: -7px; }

[dir="rtl"] .tTvXye .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .tTvXye .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc[dir="rtl"] { margin-left: -7px; margin-right: 8px; }

.tTvXye .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { margin-left: 8px; margin-right: -7px; }

[dir="rtl"] .tTvXye .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .tTvXye .VfPpkd-Zr1Nwf-OWXEXe-UbuQg[dir="rtl"] { margin-left: -7px; margin-right: 8px; }

.tTvXye .VfPpkd-v1cqY { top: -1px; left: -1px; border: 1px solid transparent; }

.tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd { padding-right: 11px; padding-left: 11px; border-width: 1px; border-color: var(--gm-chip-outline-color,rgb(232,240,254)); }

.tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus, .tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe { padding-right: 11px; padding-left: 11px; border-width: 1px; }

.tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus .VfPpkd-v1cqY, .tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe .VfPpkd-v1cqY { top: -1px; left: -1px; border: 1px solid transparent; }

.tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY { top: -1px; left: -1px; border: 1px solid transparent; }

.tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus, .tTvXye.RgtwTe.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe { border-color: var(--gm-chip-outline-color--stateful,rgb(23,78,166)); }

.KshDhe { color: var(--gm-chip-ink-color,rgb(60,64,67)); }

.KshDhe .VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { width: 20px; height: 20px; font-size: 20px; }

.KshDhe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, .KshDhe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { margin-left: -8px; margin-right: 8px; }

[dir="rtl"] .KshDhe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, [dir="rtl"] .KshDhe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce), .KshDhe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir="rtl"], .KshDhe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir="rtl"] { margin-left: 8px; margin-right: -8px; }

.KshDhe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(60, 64, 67); }

.KshDhe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color,rgb(60,64,67)); }

.KshDhe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(60, 64, 67); }

.KshDhe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(60, 64, 67); }

.KshDhe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(60, 64, 67); }

.KshDhe .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color,rgb(60,64,67)); }

.KshDhe:hover, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus, .KshDhe:active { color: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.KshDhe:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc, .KshDhe:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc { color: rgb(32, 33, 36); }

.KshDhe:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .KshDhe:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.KshDhe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg, .KshDhe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg { color: rgb(32, 33, 36); }

.KshDhe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover, .KshDhe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover { color: rgb(32, 33, 36); }

.KshDhe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus, .KshDhe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus { color: rgb(32, 33, 36); }

.KshDhe:hover .VfPpkd-PvL5qd-Jt5cK, .KshDhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK, .KshDhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK, .KshDhe:active .VfPpkd-PvL5qd-Jt5cK { stroke: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.PdGJo, .PdGJo .VfPpkd-v1cqY, .Zn20Xd, .Zn20Xd .VfPpkd-v1cqY { border-radius: 8px; }

.Zn20Xd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, .Zn20Xd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce) { margin-left: -8px; margin-right: 8px; }

[dir="rtl"] .Zn20Xd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd, [dir="rtl"] .Zn20Xd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce), .Zn20Xd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir="rtl"], .Zn20Xd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir="rtl"] { margin-left: 8px; margin-right: -8px; }

.Zx360 .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color,rgb(95,99,104)); }

.Zx360 .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .Zx360 .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { background-color: var(--gm-chip-state-color,rgb(60,64,67)); }

.Zx360:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .Zx360.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.Zx360.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before, .Zx360:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.Zx360:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { transition: opacity 0.15s linear 0s; }

.Zx360:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-XPtOyb-UbuQg-XCaCob::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.Zx360.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.Zx360:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .Zx360.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .Zx360:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc, .Zx360:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc { color: var(--gm-chip-ink-color--stateful,rgb(32,33,36)); }

.VfPpkd-StrnGf-rymPhb { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle1-font-size,1rem); font-weight: var(--mdc-typography-subtitle1-font-weight,400); letter-spacing: var(--mdc-typography-subtitle1-letter-spacing,.009375em); text-decoration: var(--mdc-typography-subtitle1-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle1-text-transform,inherit); line-height: 1.5rem; margin: 0px; padding: 8px 0px; list-style-type: none; color: var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87)); }

.VfPpkd-StrnGf-rymPhb:focus { outline: none; }

.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54)); }

.VfPpkd-StrnGf-rymPhb-f7MjDc { background-color: transparent; }

.VfPpkd-StrnGf-rymPhb-f7MjDc { color: var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38)); }

.VfPpkd-StrnGf-rymPhb-IhFlZd { color: var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38)); }

.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c { opacity: 0.38; }

.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc { padding-top: 4px; padding-bottom: 4px; font-size: 0.812rem; }

.VfPpkd-StrnGf-rymPhb-Tkg0ld { display: block; }

.VfPpkd-StrnGf-rymPhb-ibnC6b { display: flex; position: relative; -webkit-box-align: center; align-items: center; -webkit-box-pack: start; justify-content: flex-start; overflow: hidden; padding: 0px 16px; height: 48px; }

.VfPpkd-StrnGf-rymPhb-ibnC6b:focus { outline: none; }

.VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before, .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 1px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before, .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before { border-color: canvastext; }
}

.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 3px double transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before { border-color: canvastext; }
}

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 16px; padding-right: 16px; height: 56px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 16px; padding-right: 16px; height: 56px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 16px; padding-right: 16px; height: 56px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 16px; padding-right: 16px; height: 72px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 0px; padding-right: 16px; height: 72px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 20px; height: 20px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-f7MjDc { flex-shrink: 0; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; fill: currentcolor; object-fit: cover; margin-left: 0px; margin-right: 32px; width: 24px; height: 24px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 32px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 32px; width: 24px; height: 24px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 32px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 40px; height: 40px; border-radius: 50%; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 40px; height: 40px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 56px; height: 56px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 100px; height: 56px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { display: inline-flex; }

.VfPpkd-StrnGf-rymPhb-IhFlZd { margin-left: auto; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-IhFlZd:not(.HzV7m-fuEl3d) { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-caption-font-size,.75rem); line-height: var(--mdc-typography-caption-line-height,1.25rem); font-weight: var(--mdc-typography-caption-font-weight,400); letter-spacing: var(--mdc-typography-caption-letter-spacing,.0333333333em); text-decoration: var(--mdc-typography-caption-text-decoration,inherit); text-transform: var(--mdc-typography-caption-text-transform,inherit); }

.VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] .VfPpkd-StrnGf-rymPhb-IhFlZd, [dir="rtl"] .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-IhFlZd { margin-left: 0px; margin-right: auto; }

.VfPpkd-StrnGf-rymPhb-b9t22c { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; }

.VfPpkd-StrnGf-rymPhb-b9t22c[for] { pointer-events: none; }

.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 24px; content: ""; vertical-align: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-body2-font-size,.875rem); font-weight: var(--mdc-typography-body2-font-weight,400); letter-spacing: var(--mdc-typography-body2-letter-spacing,.0178571429em); text-decoration: var(--mdc-typography-body2-text-decoration,inherit); text-transform: var(--mdc-typography-body2-text-transform,inherit); text-overflow: ellipsis; white-space: nowrap; overflow: hidden; display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS::before { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { font-size: inherit; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b { height: 40px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-b9t22c { align-self: flex-start; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-ibnC6b { height: 64px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b { height: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc { align-self: flex-start; margin-top: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b { height: 60px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; width: 36px; height: 36px; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b { cursor: pointer; }

a.VfPpkd-StrnGf-rymPhb-ibnC6b { color: inherit; text-decoration: none; }

.VfPpkd-StrnGf-rymPhb-clz4Ic { height: 0px; margin: 0px; border-top: none; border-right: none; border-left: none; border-bottom: 1px solid; border-image: initial; }

.VfPpkd-StrnGf-rymPhb-clz4Ic { border-bottom-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd, .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe { margin-left: 72px; margin-right: 0px; width: calc(100% - 72px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe, .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd { margin-left: 72px; margin-right: 0px; width: calc(100% - 88px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd, .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 72px; margin-right: 0px; width: calc(100% - 72px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 72px; margin-right: 0px; width: calc(100% - 88px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 72px; margin-right: 0px; width: calc(100% - 72px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 72px; margin-right: 0px; width: calc(100% - 88px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 72px; margin-right: 0px; width: calc(100% - 72px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 72px; margin-right: 0px; width: calc(100% - 88px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 72px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 88px; margin-right: 0px; width: calc(100% - 88px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 88px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 88px; margin-right: 0px; width: calc(100% - 104px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 88px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 116px; margin-right: 0px; width: calc(100% - 116px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 116px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 116px; margin-right: 0px; width: calc(100% - 132px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 116px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 0px; margin-right: 0px; width: 100%; }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 0px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 0px; }

.VfPpkd-StrnGf-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb { padding: 0px; }

.VfPpkd-StrnGf-rymPhb-oT7voc { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle1-font-size,1rem); line-height: var(--mdc-typography-subtitle1-line-height,1.75rem); font-weight: var(--mdc-typography-subtitle1-font-weight,400); letter-spacing: var(--mdc-typography-subtitle1-letter-spacing,.009375em); text-decoration: var(--mdc-typography-subtitle1-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle1-text-transform,inherit); margin: 0.75rem 16px; }

.VfPpkd-rymPhb-fpDzbe-fmcmS { color: var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87)); }

.VfPpkd-rymPhb-L8ivfd-fmcmS { color: var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54)); }

.VfPpkd-rymPhb-bC5pod-fmcmS { color: var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38)); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e { background-color: transparent; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e { color: var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38)); }

.VfPpkd-rymPhb-JMEf7e { color: var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38)); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e { opacity: 0.38; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { color: var(--mdc-theme-on-surface,#000); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS, .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb { color: var(--mdc-theme-primary,#6200ee); }

.VfPpkd-StrnGf-rymPhb-oT7voc { color: var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87)); }

.VfPpkd-rymPhb-clz4Ic::after { border-bottom-color: white; }

.VfPpkd-rymPhb { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle1-font-size,1rem); font-weight: var(--mdc-typography-subtitle1-font-weight,400); letter-spacing: var(--mdc-typography-subtitle1-letter-spacing,.009375em); text-decoration: var(--mdc-typography-subtitle1-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle1-text-transform,inherit); line-height: 1.5rem; }

.VfPpkd-rymPhb-fpDzbe-fmcmS { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle1-font-size,1rem); line-height: var(--mdc-typography-subtitle1-line-height,1.75rem); font-weight: var(--mdc-typography-subtitle1-font-weight,400); letter-spacing: var(--mdc-typography-subtitle1-letter-spacing,.009375em); text-decoration: var(--mdc-typography-subtitle1-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle1-text-transform,inherit); }

.VfPpkd-rymPhb-L8ivfd-fmcmS { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-body2-font-size,.875rem); line-height: var(--mdc-typography-body2-line-height,1.25rem); font-weight: var(--mdc-typography-body2-font-weight,400); letter-spacing: var(--mdc-typography-body2-letter-spacing,.0178571429em); text-decoration: var(--mdc-typography-body2-text-decoration,inherit); text-transform: var(--mdc-typography-body2-text-transform,inherit); }

.VfPpkd-rymPhb-bC5pod-fmcmS { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-overline-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-overline-font-size,.75rem); line-height: var(--mdc-typography-overline-line-height,2rem); font-weight: var(--mdc-typography-overline-font-weight,500); letter-spacing: var(--mdc-typography-overline-letter-spacing,.1666666667em); text-decoration: var(--mdc-typography-overline-text-decoration,none); text-transform: var(--mdc-typography-overline-text-transform,uppercase); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb { width: 40px; height: 40px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb { width: 24px; height: 24px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb { width: 40px; height: 40px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb { width: 56px; height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb { width: 100px; height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb { width: 40px; height: 40px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb { width: 36px; height: 20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e { width: 24px; height: 24px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e { width: 40px; height: 40px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e { width: 36px; height: 20px; }

.VfPpkd-rymPhb-oT7voc { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-subtitle1-font-size,1rem); line-height: var(--mdc-typography-subtitle1-line-height,1.75rem); font-weight: var(--mdc-typography-subtitle1-font-weight,400); letter-spacing: var(--mdc-typography-subtitle1-letter-spacing,.009375em); text-decoration: var(--mdc-typography-subtitle1-text-decoration,inherit); text-transform: var(--mdc-typography-subtitle1-text-transform,inherit); }

.VfPpkd-rymPhb-clz4Ic { background-color: rgba(0, 0, 0, 0.12); }

.VfPpkd-rymPhb-clz4Ic { height: 1px; }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .VfPpkd-rymPhb-clz4Ic::after { content: ""; display: block; border-bottom-width: 1px; border-bottom-style: solid; }
}

.VfPpkd-rymPhb { margin: 0px; padding: 8px 0px; list-style-type: none; }

.VfPpkd-rymPhb:focus { outline: none; }

.VfPpkd-rymPhb-Tkg0ld { display: block; }

.VfPpkd-rymPhb-ibnC6b { display: flex; position: relative; -webkit-box-pack: start; justify-content: flex-start; overflow: hidden; padding: 0px; -webkit-box-align: stretch; align-items: stretch; cursor: pointer; }

.VfPpkd-rymPhb-ibnC6b:focus { outline: none; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 48px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 64px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb { height: 88px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-KkROqb { align-self: center; margin-top: 0px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 16px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: center; margin-top: 0px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: flex-start; margin-top: 16px; }

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me, .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-tPcied-hXIJHe { cursor: auto; }

.VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before, .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 1px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before, .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before { border-color: canvastext; }
}

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 3px double transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before { border-color: canvastext; }
}

.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 3px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before { border-color: canvastext; }
}

a.VfPpkd-rymPhb-ibnC6b { color: inherit; text-decoration: none; }

.VfPpkd-rymPhb-KkROqb { fill: currentcolor; flex-shrink: 0; pointer-events: none; }

.VfPpkd-rymPhb-JMEf7e { flex-shrink: 0; pointer-events: none; }

.VfPpkd-rymPhb-Gtdoyb { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; align-self: center; -webkit-box-flex: 1; flex: 1 1 0%; pointer-events: none; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-Gtdoyb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-Gtdoyb { align-self: stretch; }

.VfPpkd-rymPhb-Gtdoyb[for] { pointer-events: none; }

.VfPpkd-rymPhb-fpDzbe-fmcmS { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-L8ivfd-fmcmS { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-L8ivfd-fmcmS::before { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS { white-space: normal; line-height: 20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj .VfPpkd-rymPhb-L8ivfd-fmcmS { white-space: nowrap; }

.VfPpkd-rymPhb-bC5pod-fmcmS { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 24px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb { border-radius: 50%; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 32px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 32px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb { margin-left: 0px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb { margin-left: 8px; margin-right: 24px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 24px; margin-right: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb { margin-left: 8px; margin-right: 24px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 24px; margin-right: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS { display: block; margin-top: 0px; line-height: normal; margin-bottom: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: -20px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 32px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb { height: 72px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: flex-start; margin-top: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { margin-left: 28px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 16px; margin-right: 28px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e::before { display: inline-block; width: 0px; height: 28px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { -webkit-font-smoothing: antialiased; font-family: var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif)); font-size: var(--mdc-typography-caption-font-size,.75rem); line-height: var(--mdc-typography-caption-line-height,1.25rem); font-weight: var(--mdc-typography-caption-font-weight,400); letter-spacing: var(--mdc-typography-caption-letter-spacing,.0333333333em); text-decoration: var(--mdc-typography-caption-text-decoration,inherit); text-transform: var(--mdc-typography-caption-text-transform,inherit); }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e { margin-left: 24px; margin-right: 8px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 8px; margin-right: 24px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: flex-start; margin-top: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e { margin-left: 24px; margin-right: 8px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 8px; margin-right: 24px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: flex-start; margin-top: 8px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e, .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e { align-self: flex-start; margin-top: 16px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS { display: block; margin-top: 0px; line-height: normal; }

.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before { display: inline-block; width: 0px; height: 20px; content: ""; vertical-align: 0px; }

.VfPpkd-rymPhb-ibnC6b { padding-left: 16px; padding-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-ibnC6b, .VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 16px; }

.VfPpkd-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb { padding: 0px; }

.VfPpkd-rymPhb-oT7voc { margin: 0.75rem 16px; }

.VfPpkd-rymPhb-clz4Ic { padding: 0px; background-clip: content-box; }

.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe { padding-left: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"] { padding-right: 16px; }

.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe { padding-right: 16px; }

[dir="rtl"] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, [dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"], .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"] { padding-left: 16px; }

.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe { padding-left: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"] { padding-right: 0px; }

[dir="rtl"] .VfPpkd-rymPhb-clz4Ic, .VfPpkd-rymPhb-clz4Ic[dir="rtl"] { padding: 0px; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after { z-index: var(--mdc-ripple-z-index,0); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-StrnGf-rymPhb-pZXsl::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-StrnGf-rymPhb-pZXsl::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-StrnGf-rymPhb-pZXsl::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { z-index: var(--mdc-ripple-z-index,0); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after { top: -50%; left: -50%; width: 200%; height: 200%; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { top: -50%; left: -50%; width: 200%; height: 200%; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,#000); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,#000); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-activated-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.16); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.24); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.24); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-activated-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.16); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.24); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.24); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.24); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-selected-opacity,.08); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.2); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.2); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-selected-opacity,.08); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.12); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.2); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.2); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.2); }

:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl, :not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl { position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; pointer-events: none; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { z-index: var(--mdc-ripple-z-index,0); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { top: -50%; left: -50%; width: 200%; height: 200%; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,#000); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-activated-opacity,.12); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.16); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.24); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.24); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.24); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-selected-opacity,.08); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee)); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.12); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, :not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.2); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.2); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.2); }

:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl { outline: none; overflow: hidden; position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; pointer-events: none; }

.P2Hi5d, .mkMxfe, .OBi8lb, .P9QRxe, .vqjb4e, .y8Rdrf, .DMZ54e { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: var(--mdc-theme-on-surface,#000); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-IhFlZd, .mkMxfe .VfPpkd-StrnGf-rymPhb-IhFlZd, .OBi8lb .VfPpkd-StrnGf-rymPhb-IhFlZd, .P9QRxe .VfPpkd-StrnGf-rymPhb-IhFlZd, .vqjb4e .VfPpkd-StrnGf-rymPhb-IhFlZd, .y8Rdrf .VfPpkd-StrnGf-rymPhb-IhFlZd, .DMZ54e .VfPpkd-StrnGf-rymPhb-IhFlZd { color: rgb(95, 99, 104); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: rgb(60, 64, 67); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c { opacity: 0.38; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b { color: var(--mdc-theme-on-surface,#000); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc { color: var(--mdc-theme-on-surface,#000); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: 0; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd { background-color: rgb(232, 240, 254); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,rgb(26,115,232)); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: graytext; }
  .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c { opacity: 1; }
}

.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 24px; padding-right: 16px; }

[dir="rtl"] .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b, .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 24px; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 24px; margin-right: 0px; width: calc(100% - 24px); }

[dir="rtl"] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 24px; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 24px; margin-right: 0px; width: calc(100% - 40px); }

[dir="rtl"] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 24px; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 24px; margin-right: 0px; width: calc(100% - 24px); }

[dir="rtl"] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 24px; }

.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 24px; margin-right: 0px; width: calc(100% - 40px); }

[dir="rtl"] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 24px; }

.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc { margin-left: 0px; margin-right: 16px; }

[dir="rtl"] .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc, .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir="rtl"] { margin-left: 16px; margin-right: 0px; }

.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc { margin-left: 56px; margin-right: 0px; width: calc(100% - 56px); }

[dir="rtl"] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc, .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir="rtl"] { margin-left: 0px; margin-right: 56px; }

.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { width: calc(100% - 16px); }

.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg { margin-left: 56px; margin-right: 0px; width: calc(100% - 72px); }

[dir="rtl"] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg, .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir="rtl"] { margin-left: 0px; margin-right: 56px; }

.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 16px); }

[dir="rtl"] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2, .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2 { margin-left: 16px; margin-right: 0px; width: calc(100% - 32px); }

[dir="rtl"] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2, .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir="rtl"] { margin-left: 0px; margin-right: 16px; }

.r6B9Fd { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; }

.r6B9Fd .VfPpkd-rymPhb-fpDzbe-fmcmS { color: rgb(60, 64, 67); }

.r6B9Fd .VfPpkd-rymPhb-L8ivfd-fmcmS, .r6B9Fd .VfPpkd-rymPhb-bC5pod-fmcmS, .r6B9Fd .VfPpkd-rymPhb-JMEf7e { color: rgb(95, 99, 104); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { color: rgb(60, 64, 67); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e { opacity: 0.38; }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb { color: rgb(60, 64, 67); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before { opacity: 0; }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd { background-color: rgb(232, 240, 254); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before, .r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,rgb(26,115,232)); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before, .r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before, .r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

@media screen and (forced-colors: active) {
  .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e { color: graytext; }
  .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb, .r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e { opacity: 1; }
}

.uTZ9Lb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb, .FvXOfd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb, .QrsYgb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb, .gfwIBd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: center; margin-top: 0px; }

.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 56px; }

.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc, .HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc { height: 72px; }

.UbEQCe.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .UbEQCe.VfPpkd-rymPhb-ibnC6b, .UbEQCe.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.UbEQCe .VfPpkd-rymPhb-KkROqb { margin-left: 16px; margin-right: 16px; }

[dir="rtl"] .UbEQCe .VfPpkd-rymPhb-KkROqb, .UbEQCe .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 16px; margin-right: 16px; }

.rKASPc.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .rKASPc.VfPpkd-rymPhb-ibnC6b, .rKASPc.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.rKASPc .VfPpkd-rymPhb-KkROqb { margin-left: 8px; margin-right: 8px; }

[dir="rtl"] .rKASPc .VfPpkd-rymPhb-KkROqb, .rKASPc .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 8px; margin-right: 8px; }

.rKASPc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.U5k4Fd.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .U5k4Fd.VfPpkd-rymPhb-ibnC6b, .U5k4Fd.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.U5k4Fd .VfPpkd-rymPhb-KkROqb { margin-left: 8px; margin-right: 8px; }

[dir="rtl"] .U5k4Fd .VfPpkd-rymPhb-KkROqb, .U5k4Fd .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 8px; margin-right: 8px; }

.U5k4Fd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.ifEyr.VfPpkd-rymPhb-ibnC6b { padding-left: 0px; }

[dir="rtl"] .ifEyr.VfPpkd-rymPhb-ibnC6b, .ifEyr.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-right: 0px; }

.ifEyr .VfPpkd-rymPhb-KkROqb { margin-left: 8px; margin-right: 8px; }

[dir="rtl"] .ifEyr .VfPpkd-rymPhb-KkROqb, .ifEyr .VfPpkd-rymPhb-KkROqb[dir="rtl"] { margin-left: 8px; margin-right: 8px; }

.ifEyr.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb { align-self: flex-start; margin-top: 8px; }

.SNowt.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .SNowt.VfPpkd-rymPhb-ibnC6b, .SNowt.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.SNowt .VfPpkd-rymPhb-JMEf7e { margin-left: 8px; margin-right: 16px; }

[dir="rtl"] .SNowt .VfPpkd-rymPhb-JMEf7e, .SNowt .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 16px; margin-right: 8px; }

.tfmWAf.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .tfmWAf.VfPpkd-rymPhb-ibnC6b, .tfmWAf.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.tfmWAf .VfPpkd-rymPhb-JMEf7e { margin-left: 8px; margin-right: 16px; }

[dir="rtl"] .tfmWAf .VfPpkd-rymPhb-JMEf7e, .tfmWAf .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 16px; margin-right: 8px; }

.axtYbd.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .axtYbd.VfPpkd-rymPhb-ibnC6b, .axtYbd.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.axtYbd .VfPpkd-rymPhb-JMEf7e { margin-left: 16px; margin-right: 24px; }

[dir="rtl"] .axtYbd .VfPpkd-rymPhb-JMEf7e, .axtYbd .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 24px; margin-right: 16px; }

.aopLEb.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .aopLEb.VfPpkd-rymPhb-ibnC6b, .aopLEb.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.aopLEb .VfPpkd-rymPhb-JMEf7e { margin-left: 16px; margin-right: 24px; }

[dir="rtl"] .aopLEb .VfPpkd-rymPhb-JMEf7e, .aopLEb .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 24px; margin-right: 16px; }

.zlqiud.VfPpkd-rymPhb-ibnC6b { padding-right: 0px; }

[dir="rtl"] .zlqiud.VfPpkd-rymPhb-ibnC6b, .zlqiud.VfPpkd-rymPhb-ibnC6b[dir="rtl"] { padding-left: 0px; }

.zlqiud .VfPpkd-rymPhb-JMEf7e { margin-left: 16px; margin-right: 24px; }

[dir="rtl"] .zlqiud .VfPpkd-rymPhb-JMEf7e, .zlqiud .VfPpkd-rymPhb-JMEf7e[dir="rtl"] { margin-left: 24px; margin-right: 16px; }

.isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe { padding-left: 24px; }

[dir="rtl"] .isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe, .isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir="rtl"] { padding-right: 24px; }

.MCs1Pd { padding-left: 24px; padding-right: 24px; }

[dir="rtl"] .MCs1Pd, .MCs1Pd[dir="rtl"] { padding-left: 24px; padding-right: 24px; }

.e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe { padding-right: 24px; }

[dir="rtl"] .e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe, .e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir="rtl"] { padding-left: 24px; }

[dir="rtl"] .e6pQl, .e6pQl[dir="rtl"] { padding: 0px; }

.VfPpkd-xl07Ob-XxIAqe { display: none; position: absolute; box-sizing: border-box; margin: 0px; padding: 0px; transform: scale(1); transform-origin: left top; opacity: 0; overflow: auto; will-change: transform, opacity; box-shadow: rgba(0, 0, 0, 0.2) 0px 5px 5px -3px, rgba(0, 0, 0, 0.14) 0px 8px 10px 1px, rgba(0, 0, 0, 0.12) 0px 3px 14px 2px; }

.VfPpkd-xl07Ob-XxIAqe:focus { outline: none; }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-FNFY6c { display: inline-block; transform: scale(0.8); opacity: 0; }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-FNFY6c { display: inline-block; transform: scale(1); opacity: 1; }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO { display: inline-block; opacity: 0; }

[dir="rtl"] .VfPpkd-xl07Ob-XxIAqe, .VfPpkd-xl07Ob-XxIAqe[dir="rtl"] { }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd { position: relative; overflow: visible; }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL { position: fixed; }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-tsQazb { width: 100%; }

.VfPpkd-xl07Ob-XxIAqe { max-width: var(--mdc-menu-max-width,calc(100vw - 32px)); max-height: var(--mdc-menu-max-height,calc(100vh - 32px)); z-index: 8; transition: opacity 0.03s linear 0s, transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0s, height 0.25s cubic-bezier(0, 0, 0.2, 1) 0s, -webkit-transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0s; background-color: var(--mdc-theme-surface,#fff); color: var(--mdc-theme-on-surface,#000); border-radius: var(--mdc-shape-medium,4px); }

.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO { transition: opacity 75ms linear 0s; }

.UQ5E0 { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 5px -1px, rgba(0, 0, 0, 0.14) 0px 6px 10px 0px, rgba(0, 0, 0, 0.12) 0px 1px 18px 0px; }

.VfPpkd-xl07Ob { min-width: var(--mdc-menu-min-width,112px); }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-IhFlZd, .VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-f7MjDc { color: rgba(0, 0, 0, 0.87); }

.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: 0.04; }

.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-rymPhb-pZXsl::before { opacity: 0.04; }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb { color: rgba(0, 0, 0, 0.87); }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb, .VfPpkd-xl07Ob .VfPpkd-rymPhb { position: relative; }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb, .VfPpkd-xl07Ob .VfPpkd-rymPhb .VfPpkd-BFbNVe-bF1uUb { width: 100%; height: 100%; top: 0px; left: 0px; }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before, .VfPpkd-xl07Ob .VfPpkd-rymPhb::before { position: absolute; box-sizing: border-box; width: 100%; height: 100%; top: 0px; left: 0px; border: 1px solid transparent; border-radius: inherit; content: ""; pointer-events: none; }

@media screen and (forced-colors: active) {
  .VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before, .VfPpkd-xl07Ob .VfPpkd-rymPhb::before { border-color: canvastext; }
}

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-clz4Ic { margin: 8px 0px; }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b { user-select: none; }

.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me { cursor: auto; }

.VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-b9t22c, .VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc { pointer-events: none; }

.VfPpkd-qPzbhe-JNdkSc { padding: 0px; fill: currentcolor; }

.VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b { padding-left: 56px; padding-right: 16px; }

[dir="rtl"] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b, .VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b[dir="rtl"] { padding-left: 16px; padding-right: 56px; }

.VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c { left: 16px; right: auto; visibility: hidden; position: absolute; top: 50%; transform: translateY(-50%); transition-property: visibility; transition-delay: 75ms; }

[dir="rtl"] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c, .VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c[dir="rtl"] { left: auto; right: 16px; }

.VfPpkd-xl07Ob-ibnC6b-OWXEXe-gk6SMd .VfPpkd-qPzbhe-JNdkSc-Bz112c { display: inline; visibility: visible; }

.q6oraf { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 5px -1px, rgba(0, 0, 0, 0.14) 0px 6px 10px 0px, rgba(0, 0, 0, 0.12) 0px 1px 18px 0px; }

.q6oraf .VfPpkd-StrnGf-rymPhb { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: var(--mdc-theme-on-surface,#000); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd { color: rgb(95, 99, 104); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: rgb(60, 64, 67); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c { opacity: 0.38; }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b { color: var(--mdc-theme-on-surface,#000); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc { color: var(--mdc-theme-on-surface,#000); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: 0; }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd { background-color: rgb(232, 240, 254); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after { background-color: var(--mdc-ripple-color,rgb(26,115,232)); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition: opacity 0.15s linear 0s; }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: graytext; }
  .q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c { opacity: 1; }
}

.Qo4GQ { cursor: text; position: relative; }

.NtoL8e { width: 100%; }

.FCIEcc { overflow-x: hidden; width: inherit; }

.opjjDf { padding: 0px; }

.opjjDf.fO0tQe { margin: 4px 0px 4px -0.25em; }

.opjjDf.fO0tQe .wp9Phd { padding-left: 0.25em; }

.opjjDf.fO0tQe .wp9Phd.aPRBcb { margin-left: -9px; padding-left: 0px; }

.FCIEcc .Zwu5hc.VfPpkd-StrnGf-rymPhb-f7MjDc { margin-right: 16px; width: 40px; }

.O2hkRb { position: absolute; top: -1000px; height: 1px; overflow: hidden; }

.fhj04 { -webkit-box-align: center; align-items: center; display: flex; }

.vhoiae .FCIEcc .VfPpkd-StrnGf-rymPhb, .X9XeLb .FCIEcc .VfPpkd-StrnGf-rymPhb, .cWKK1c .FCIEcc .VfPpkd-StrnGf-rymPhb, .aJfoSc .FCIEcc .VfPpkd-StrnGf-rymPhb, .TOb6Ze .FCIEcc .VfPpkd-StrnGf-rymPhb { background: var(--dt-surface3,#fff); }

.vhoiae .FCIEcc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .X9XeLb .FCIEcc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .cWKK1c .FCIEcc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .aJfoSc .FCIEcc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS, .TOb6Ze .FCIEcc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS { color: var(--dt-on-surface,rgb(60,64,67)); }

.vhoiae .FCIEcc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .X9XeLb .FCIEcc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .cWKK1c .FCIEcc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .aJfoSc .FCIEcc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS, .TOb6Ze .FCIEcc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.m0PB1.m0PB1 { background-color: var(--dt-surface1,#fff); max-width: calc(100% - 1px); border-color: var(--dt-outline,rgb(128,134,139)); padding-left: 11px; padding-right: 11px; }

.m0PB1.m0PB1:focus-within { background-color: var(--dt-secondary-container,rgb(241,243,244)); border-color: var(--dt-primary-action-stateful,rgb(24,90,188)); color: var(--dt-on-secondary-container,rgb(60,64,67)); }

.m0PB1.m0PB1:focus-within .Zx360 { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.m0PB1.m0PB1:hover .Zx360 { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.m0PB1.m0PB1 .Zx360, .m0PB1.m0PB1 .VfPpkd-TfeOUb { color: var(--dt-on-surface-variant,rgb(95,99,104)); }

.m0PB1.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe { outline: transparent solid 1px; }

.m0PB1.KZKcRc { padding-left: 1px; }

.m0PB1.KZKcRc.DgLpub { padding-left: 8px; }

.RKcto { display: flex; }

.KTPIlc { border-radius: 10px; margin-left: -4px; margin-right: 4px; height: 20px; width: 20px; }

.m0PB1.KZKcRc .KTPIlc { border-radius: 14px; margin-left: 0px; height: 28px; width: 28px; }

.m0PB1 .KTPIlc.rNe0id { border-radius: 0px; color: rgb(251, 188, 4); width: 24px; }

.m0PB1.DgLpub .KTPIlc.rNe0id { color: var(--dt-error,rgb(217,48,37)); }

.KTPIlc.PMBZAf { height: 20px; width: 20px; }

@media (forced-colors: active) {
  .m0PB1 .Zx360 { color: buttontext; }
  .m0PB1:hover .Zx360 { color: buttontext; }
  .m0PB1 .Zx360:hover, .m0PB1 .Zx360:focus { background: highlight; border: 1px solid highlighttext; color: highlighttext; }
}

.PMBZAf .co39ub { border-color: rgb(66, 133, 244); }

.PMBZAf .Cn087 { border-color: rgb(251, 188, 4); }

.PMBZAf .hfsr6b { border-color: rgb(234, 67, 53); }

.PMBZAf .EjXFBf { border-color: rgb(52, 168, 83); }

.NMm5M { fill: currentcolor; flex-shrink: 0; }

html[dir="rtl"] .hhikbc { transform: scaleX(-1); }

.EmVfjc { display: inline-block; position: relative; width: 28px; height: 28px; }

.Cg7hO { position: absolute; width: 0px; height: 0px; overflow: hidden; }

.xu46lf { width: 100%; height: 100%; }

.EmVfjc.qs41qe .xu46lf { animation: 1568ms linear 0s infinite normal none running spinner-container-rotate; }

.ir3uv { position: absolute; width: 100%; height: 100%; opacity: 0; }

.uWlRce { border-color: rgb(66, 133, 244); }

.GFoASc { border-color: rgb(219, 68, 55); }

.WpeOqd { border-color: rgb(244, 180, 0); }

.rHV3jf { border-color: rgb(15, 157, 88); }

.EmVfjc.qs41qe .ir3uv.uWlRce { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-blue-fade-in-out; }

.EmVfjc.qs41qe .ir3uv.GFoASc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-red-fade-in-out; }

.EmVfjc.qs41qe .ir3uv.WpeOqd { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-yellow-fade-in-out; }

.EmVfjc.qs41qe .ir3uv.rHV3jf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-green-fade-in-out; }

.HBnAAc { position: absolute; box-sizing: border-box; top: 0px; left: 45%; width: 10%; height: 100%; overflow: hidden; border-color: inherit; }

.HBnAAc .X6jHbb { width: 1000%; left: -450%; }

.xq3j6 { display: inline-block; position: relative; width: 50%; height: 100%; overflow: hidden; border-color: inherit; }

.xq3j6 .X6jHbb { width: 200%; }

.X6jHbb { position: absolute; inset: 0px; box-sizing: border-box; height: 100%; border-width: 3px; border-style: solid; border-top-color: inherit; border-right-color: inherit; border-left-color: inherit; border-bottom-color: transparent; border-radius: 50%; animation: 0s ease 0s 1 normal none running none; }

.xq3j6.ERcjC .X6jHbb { border-right-color: transparent; transform: rotate(129deg); }

.xq3j6.dj3yTd .X6jHbb { left: -100%; border-left-color: transparent; transform: rotate(-129deg); }

.EmVfjc.qs41qe .xq3j6.ERcjC .X6jHbb { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-left-spin; }

.EmVfjc.qs41qe .xq3j6.dj3yTd .X6jHbb { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running spinner-right-spin; }

.EmVfjc.sf4e6b .xu46lf { animation: 1568ms linear 0s infinite normal none running spinner-container-rotate, 400ms cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running spinner-fade-out; }

@-webkit-keyframes spinner-container-rotate { 
  100% { transform: rotate(360deg); }
}

@keyframes spinner-container-rotate { 
  100% { transform: rotate(360deg); }
}

@-webkit-keyframes spinner-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@keyframes spinner-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@-webkit-keyframes spinner-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@keyframes spinner-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@-webkit-keyframes spinner-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@keyframes spinner-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@-webkit-keyframes spinner-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@keyframes spinner-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@-webkit-keyframes spinner-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes spinner-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@-webkit-keyframes spinner-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@keyframes spinner-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@-webkit-keyframes spinner-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@keyframes spinner-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@-webkit-keyframes spinner-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes spinner-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

.VfPpkd-GCYh9b { padding: 10px; }

.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: rgba(0, 0, 0, 0.54); }

.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--mdc-theme-secondary,#018786); }

.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: var(--mdc-theme-secondary,#018786); }

.VfPpkd-GCYh9b [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: rgba(0, 0, 0, 0.38); }

.VfPpkd-GCYh9b [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: rgba(0, 0, 0, 0.38); }

.VfPpkd-GCYh9b [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: rgba(0, 0, 0, 0.38); }

.VfPpkd-GCYh9b .VfPpkd-RsCWK::before { background-color: var(--mdc-theme-secondary,#018786); }

.VfPpkd-GCYh9b .VfPpkd-RsCWK::before { top: -10px; left: -10px; width: 40px; height: 40px; }

.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe { top: 0px; right: 0px; left: 0px; width: 40px; height: 40px; }

@media (-ms-high-contrast:active), screen and (forced-colors: active) {
  .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: graytext; }
  .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: graytext; }
  .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: graytext; }
}

.VfPpkd-GCYh9b { display: inline-block; position: relative; -webkit-box-flex: 0; flex: 0 0 auto; box-sizing: content-box; width: 20px; height: 20px; cursor: pointer; will-change: opacity, transform, border-color, color; }

.VfPpkd-GCYh9b[hidden] { display: none; }

.VfPpkd-RsCWK { display: inline-block; position: relative; box-sizing: border-box; width: 20px; height: 20px; }

.VfPpkd-RsCWK::before { position: absolute; transform: scale(0, 0); border-radius: 50%; opacity: 0; pointer-events: none; content: ""; transition: opacity 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms, transform 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-wVo5xe-LkdAo { position: absolute; top: 0px; left: 0px; box-sizing: border-box; width: 100%; height: 100%; border-width: 2px; border-style: solid; border-radius: 50%; transition: border-color 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-Z5TpLc-LkdAo { position: absolute; top: 0px; left: 0px; box-sizing: border-box; width: 100%; height: 100%; transform: scale(0, 0); border-width: 10px; border-style: solid; border-radius: 50%; transition: transform 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms, border-color 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0.4, 0, 0.6, 1) 0ms; }

.VfPpkd-gBXA9-bMcfAe { position: absolute; margin: 0px; padding: 0px; opacity: 0; cursor: inherit; z-index: 1; }

.VfPpkd-GCYh9b-OWXEXe-dgl2Hf { margin: 4px; }

.VfPpkd-GCYh9b-OWXEXe-dgl2Hf .VfPpkd-gBXA9-bMcfAe { top: -4px; right: -4px; left: -4px; width: 48px; height: 48px; }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec, .VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec { pointer-events: none; border: 2px solid transparent; border-radius: 6px; box-sizing: content-box; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: 100%; width: 100%; }

@media screen and (forced-colors: active) {
  .VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec, .VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec { border-color: canvastext; }
}

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec::after, .VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec::after { content: ""; border: 2px solid transparent; border-radius: 8px; display: block; position: absolute; top: 50%; left: 50%; transform: translate(-50%, -50%); height: calc(100% + 4px); width: calc(100% + 4px); }

@media screen and (forced-colors: active) {
  .VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec::after, .VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec::after { border-color: canvastext; }
}

.VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK, .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK { transition: opacity 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { transition: border-color 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { transition: transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, border-color 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-GCYh9b-OWXEXe-OWB6Me { cursor: default; pointer-events: none; }

.VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { transform: scale(0.5); transition: transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, border-color 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK, [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe + .VfPpkd-RsCWK { cursor: default; }

.VfPpkd-gBXA9-bMcfAe:focus + .VfPpkd-RsCWK::before { transform: scale(1); opacity: 0.12; transition: opacity 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms, -webkit-transform 0.12s cubic-bezier(0, 0, 0.2, 1) 0ms; }

.VfPpkd-GCYh9b { --mdc-ripple-fg-size: 0; --mdc-ripple-left: 0; --mdc-ripple-top: 0; --mdc-ripple-fg-scale: 1; --mdc-ripple-fg-translate-end: 0; --mdc-ripple-fg-translate-start: 0; -webkit-tap-highlight-color: rgba(0, 0, 0, 0); will-change: transform, opacity; }

.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b .VfPpkd-eHTEvd::after { position: absolute; border-radius: 50%; opacity: 0; pointer-events: none; content: ""; }

.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before { transition: opacity 15ms linear 0s, background-color 15ms linear 0s; z-index: var(--mdc-ripple-z-index,1); }

.VfPpkd-GCYh9b .VfPpkd-eHTEvd::after { z-index: var(--mdc-ripple-z-index,0); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::before { transform: scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after { top: 0px; left: 0px; transform: scale(0); transform-origin: center center; }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-eHTEvd::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-eHTEvd::after { animation: 225ms ease 0s 1 normal forwards running mdc-ripple-fg-radius-in, 75ms ease 0s 1 normal forwards running mdc-ripple-fg-opacity-in; }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-eHTEvd::after { animation: 0.15s ease 0s 1 normal none running mdc-ripple-fg-opacity-out; transform: translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1)); }

.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b .VfPpkd-eHTEvd::after { top: 0px; left: 0px; width: 100%; height: 100%; }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after { top: var(--mdc-ripple-top,0); left: var(--mdc-ripple-left,0); width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after { width: var(--mdc-ripple-fg-size,100%); height: var(--mdc-ripple-fg-size,100%); }

.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b .VfPpkd-eHTEvd::after { background-color: var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786)); }

.VfPpkd-GCYh9b:hover .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-eHTEvd::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before, .VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-eHTEvd::after { transition: opacity 0.15s linear 0s; }

.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-eHTEvd::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.12); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.12); }

.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-RsCWK::before, .VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-RsCWK::before { content: none; }

.VfPpkd-eHTEvd { position: absolute; top: 0px; left: 0px; width: 100%; height: 100%; pointer-events: none; }

.kDzhGf { z-index: 0; }

.kDzhGf .VfPpkd-eHTEvd::before, .kDzhGf .VfPpkd-eHTEvd::after { z-index: -1; }

.kDzhGf .VfPpkd-eHTEvd::before, .kDzhGf .VfPpkd-eHTEvd::after { background-color: var(--gm-radio-state-color,rgb(26,115,232)); }

.kDzhGf:hover .VfPpkd-eHTEvd::before, .kDzhGf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-eHTEvd::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before, .kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-eHTEvd::after { transition: opacity 0.15s linear 0s; }

.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-eHTEvd::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::before, .kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::after { background-color: var(--gm-radio-state-color,rgb(60,64,67)); }

.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::before, .kDzhGf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::before { opacity: var(--mdc-ripple-hover-opacity,.04); }

.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::before, .kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::before { transition-duration: 75ms; opacity: var(--mdc-ripple-focus-opacity,.12); }

.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::after { transition: opacity 0.15s linear 0s; }

.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) ~ .VfPpkd-eHTEvd::after { transition-duration: 75ms; opacity: var(--mdc-ripple-press-opacity,.1); }

.kDzhGf.VfPpkd-ksKsZd-mWPk3d { --mdc-ripple-fg-opacity: var(--mdc-ripple-press-opacity,0.1); }

.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-stroke-color--unchecked,rgb(95,99,104)); }

.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-stroke-color--checked,rgb(26,115,232)); }

.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: var(--gm-radio-ink-color,rgb(26,115,232)); }

.kDzhGf [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-disabled-stroke-color--unchecked,rgba(60,64,67,.38)); }

.kDzhGf [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-disabled-stroke-color--checked,rgba(60,64,67,.38)); }

.kDzhGf [aria-disabled="true"] .VfPpkd-gBXA9-bMcfAe + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: var(--gm-radio-disabled-ink-color,rgba(60,64,67,.38)); }

.kDzhGf .VfPpkd-RsCWK::before { background-color: var(--gm-radio-state-color,rgb(26,115,232)); }

.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked) + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-stroke-color--unchecked-stateful,rgb(32,33,36)); }

.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo, .kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled:checked + .VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo { border-color: var(--gm-radio-stroke-color--checked-stateful,rgb(23,78,166)); }

.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo, .kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled + .VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo { border-color: var(--gm-radio-ink-color--stateful,rgb(23,78,166)); }

.wHsUjf { will-change: unset; }

.As7zrc { box-sizing: border-box; display: inline-flex; max-width: 100%; }

.As7zrc.UMYKE { flex-wrap: wrap; }

.SLLE9e { --mdc-checkbox-unselected-icon-color: var(--dt-on-surface-variant,rgb(95,99,104)); --mdc-checkbox-unselected-hover-icon-color: var(--dt-on-surface,rgb(60,64,67)); --mdc-checkbox-unselected-focus-icon-color: var(--dt-on-surface,rgb(60,64,67)); --mdc-checkbox-selected-checkmark-color: var(--dt-background,#fff); --mdc-checkbox-selected-icon-color: var(--dt-primary-action,rgb(25,103,210)); --mdc-checkbox-selected-hover-icon-color: var(--dt-primary-action-stateful,rgb(24,90,188)); --mdc-checkbox-selected-focus-icon-color: var(--dt-primary-action-stateful,rgb(24,90,188)); --mdc-checkbox-unselected-pressed-icon-color: var(--dt-on-surface,rgb(60,64,67)); --mdc-checkbox-selected-pressed-icon-color: var(--dt-primary-action-stateful,rgb(24,90,188)); --mdc-checkbox-disabled-unselected-icon-color: var(--dt-on-disabled,rgba(60,64,67,0.38)); --mdc-checkbox-disabled-selected-icon-color: var(--dt-on-disabled,rgba(60,64,67,0.38)); --mdc-checkbox-unselected-hover-state-layer-color: var(--dt-on-surface,rgb(60,64,67)); --mdc-checkbox-selected-hover-state-layer-color: var(--dt-primary-action,rgb(25,103,210)); --mdc-ripple-color: var(--dt-on-surface,rgb(60,64,67)); --gm-radio-state-color: var(--dt-primary-action-stateful,rgb(24,90,188)); --gm-radio-ink-color: var(--dt-primary-action,rgb(25,103,210)); --gm-radio-ink-color--stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); --gm-radio-stroke-color--checked: var(--dt-primary-action,rgb(25,103,210)); --gm-radio-stroke-color--checked-stateful: var(--dt-primary-action-stateful,rgb(24,90,188)); --gm-radio-stroke-color--unchecked: var(--dt-on-surface-variant,rgb(95,99,104)); --gm-radio-stroke-color--unchecked-stateful: var(--dt-on-surface,rgb(60,64,67)); --gm-radio-disabled-ink-color: var(--dt-on-disabled,rgba(60,64,67,0.38)); --gm-radio-disabled-stroke-color--checked: var(--dt-on-disabled,rgba(60,64,67,0.38)); --gm-radio-disabled-stroke-color--unchecked: var(--dt-on-disabled,rgba(60,64,67,0.38)); }

.SLLE9e.NWlIHc { padding: calc((var(--mdc-checkbox-ripple-size, 36px) - 18px)/2); margin: calc((var(--mdc-checkbox-touch-target-size, 36px) - 36px)/2); }

.SLLE9e.NWlIHc .VfPpkd-YQoJzd { top: calc((var(--mdc-checkbox-ripple-size, 36px) - 18px)/2); left: calc((var(--mdc-checkbox-ripple-size, 36px) - 18px)/2); }

.SLLE9e.NWlIHc .VfPpkd-muHVFf-bMcfAe { top: calc((36px - var(--mdc-checkbox-touch-target-size, 36px))/2); right: calc((36px - var(--mdc-checkbox-touch-target-size, 36px))/2); left: calc((36px - var(--mdc-checkbox-touch-target-size, 36px))/2); width: var(--mdc-checkbox-touch-target-size,36px); height: var(--mdc-checkbox-touch-target-size,36px); }

.SLLE9e.nsKVp { padding: calc((var(--mdc-checkbox-ripple-size, 32px) - 18px)/2); margin: calc((var(--mdc-checkbox-touch-target-size, 32px) - 32px)/2); }

.SLLE9e.nsKVp .VfPpkd-YQoJzd { top: calc((var(--mdc-checkbox-ripple-size, 32px) - 18px)/2); left: calc((var(--mdc-checkbox-ripple-size, 32px) - 18px)/2); }

.SLLE9e.nsKVp .VfPpkd-muHVFf-bMcfAe { top: calc((32px - var(--mdc-checkbox-touch-target-size, 32px))/2); right: calc((32px - var(--mdc-checkbox-touch-target-size, 32px))/2); left: calc((32px - var(--mdc-checkbox-touch-target-size, 32px))/2); width: var(--mdc-checkbox-touch-target-size,32px); height: var(--mdc-checkbox-touch-target-size,32px); }

.SLLE9e.GND07b { padding: calc((var(--mdc-checkbox-ripple-size, 28px) - 18px)/2); margin: calc((var(--mdc-checkbox-touch-target-size, 28px) - 28px)/2); }

.SLLE9e.GND07b .VfPpkd-YQoJzd { top: calc((var(--mdc-checkbox-ripple-size, 28px) - 18px)/2); left: calc((var(--mdc-checkbox-ripple-size, 28px) - 18px)/2); }

.SLLE9e.GND07b .VfPpkd-muHVFf-bMcfAe { top: calc((28px - var(--mdc-checkbox-touch-target-size, 28px))/2); right: calc((28px - var(--mdc-checkbox-touch-target-size, 28px))/2); left: calc((28px - var(--mdc-checkbox-touch-target-size, 28px))/2); width: var(--mdc-checkbox-touch-target-size,28px); height: var(--mdc-checkbox-touch-target-size,28px); }

.fbtU2b { font: var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-medium-spacing,.0142857143em); color: var(--dt-on-surface,rgb(60,64,67)); }

.fbtU2b:not(.RDPZE) [checkbox-label] { cursor: pointer; }

.fbtU2b.RDPZE.vf9sSe { color: var(--dt-on-disabled,rgba(60,64,67,.38)); }

.JehjSc { -webkit-box-flex: 0; flex: 0 0 100%; height: 0px; }

.EpkZi { font: var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif; letter-spacing: var(--dt-body-small-spacing,.025em); color: var(--dt-on-surface-variant,rgb(95,99,104)); margin: 0px; padding-left: 52px; position: relative; top: -10px; }

.EpkZi.gjjPnc { padding-left: 0px; }

.C0oVfc { line-height: 20px; min-width: 88px; }

.C0oVfc .RveJvd { margin: 8px; }

.fb0g6 { position: relative; }

.HB1eCd-UMrnmb .HB1eCd-UMrnmb-PvRhvb-Bz112c { display: flex; align-items: center; margin-right: 12px; height: 24px; width: 24px; }

.HB1eCd-UMrnmb .HB1eCd-UMrnmb-PvRhvb-Bz112c .HB1eCd-UMrnmb-PvRhvb-Bz112c-r9oPif { height: 24px; margin: 0px; width: 24px; }

.HB1eCd-UMrnmb .HB1eCd-UMrnmb-PvRhvb-Bz112c-Jt5cK { fill: rgb(26, 115, 232); }

.uN1Vpe { width: 520px; max-height: 90vh; overflow: auto; background-color: rgb(255, 255, 255); position: fixed; z-index: 10001; border-radius: 8px; outline: none; box-shadow: rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 3px 1px -2px, rgba(0, 0, 0, 0.2) 0px 1px 5px 0px; }

.U7DqAf { display: flex; align-items: center; justify-content: center; position: fixed; inset: 0px; background-color: rgba(0, 0, 0, 0.54); z-index: 10000; }

.Ryuoke { position: absolute; top: 16px; right: 16px; cursor: pointer; background-image: url("https://www.gstatic.com/images/icons/material/system/2x/close_grey600_24dp.png"); background-size: 24px; background-repeat: no-repeat; border: none; background-color: transparent; text-indent: -20000vh; width: 24px; height: 24px; }

.OUJMYd { flex-direction: column; display: flex; padding: 24px; font-size: 16px; color: rgb(60, 64, 67); }

.e5m6Fd { font-family: "Google Sans", sans-serif; font-size: 22px; line-height: 28px; color: rgb(32, 33, 36); margin-bottom: 16px; }

.OrGqHe { font-style: italic; margin-bottom: 12px; }

.NMjLRd { display: flex; flex-direction: row; margin: 12px 0px; }

.fhwvPe { flex: 0 0 auto; margin: 4px 0px; }

.j3YOB { flex: 1 1 auto; margin-left: 8px; cursor: pointer; }

.BeGV9d { margin-bottom: 16px; }

.G6Bwjd { border-radius: 4px; border: 1px solid rgb(218, 220, 224); box-sizing: border-box; height: 120px; padding: 8px; width: 100%; }

.msk02b { padding-bottom: 12px; }

.G6Bwjd:focus::placeholder { color: transparent; }

.G6Bwjd::placeholder { color: rgb(95, 99, 104); font-size: 16px; line-height: 30px; text-indent: 12px; }

.Ctrb4 { margin-bottom: 16px; }

.uvJjEb { display: flex; flex-direction: row; }

.m53shd { flex: 0 0 auto; margin: 4px 0px; }

.nyOE7 { flex: 1 1 auto; margin-left: 8px; }

.Aq1eFf { cursor: pointer; display: block; margin-bottom: 8px; }

.V3FtHb { color: rgb(128, 134, 139); font-size: 12px; line-height: 16px; margin-bottom: 8px; }

.iknmdd { font-size: 12px; font-weight: 500; line-height: 16px; color: rgb(197, 34, 31); margin-bottom: 8px; }

.SlYZf { color: rgb(26, 115, 232); text-decoration: underline; font-size: 12px; display: none; }

.rYRXsc { border: 1px solid lightgray; padding: 8px; max-height: 200px; overflow: auto; display: none; }

.uvJjEb.N2RpBe .Fpf1ub { display: inline; }

.uvJjEb.N2RpBe.qc48ac .Fpf1ub { display: none; }

.uvJjEb.N2RpBe.qc48ac .oeFy3e { display: inline; }

.uvJjEb.N2RpBe.qc48ac ~ .rYRXsc { display: block; }

.vAiHcc { display: flex; flex-direction: row; justify-content: flex-end; }

.jbJh6c { padding: 8px 20px; margin-left: 10px; border: none; border-radius: 4px; font: 500 14px / 20px "Google Sans", sans-serif; text-decoration: none; cursor: pointer; outline: none; }

.jbJh6c.LX7cvc { color: rgb(95, 99, 104); background-color: rgb(255, 255, 255); }

.jbJh6c.LX7cvc:hover, .jbJh6c.LX7cvc:focus { background: rgb(245, 245, 245); }

.jbJh6c.LX7cvc:active { background: rgb(214, 214, 214); }

.jbJh6c.tL9Jbf { color: rgb(255, 255, 255); background-color: rgb(26, 115, 232); }

.jbJh6c.tL9Jbf:hover, .jbJh6c.tL9Jbf:focus { background: rgb(43, 125, 233); box-shadow: rgb(223, 233, 250) 0px 1px 3px 1px; }

.jbJh6c.tL9Jbf:active { background: rgb(99, 160, 239); box-shadow: rgb(223, 233, 250) 0px 2px 6px 2px; }

.jbJh6c.tL9Jbf:disabled { background-color: rgb(189, 193, 198); }

.qb7Peb { text-rendering: geometricprecision; color: rgb(32, 33, 36); border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 2px 0px, rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; background-color: rgb(255, 255, 255); position: relative; z-index: 10000; }

.KS1ex { height: 100%; display: inline-block; outline: none; }

.dHgrtd { display: flex; flex-wrap: nowrap; padding: 4px 6px; }

.EXTU7, .UuUQYe { cursor: pointer; line-height: 18px; padding: 4px; }

.EXTU7 { border-radius: 4px; }

.EXTU7:hover, .UuUQYe:hover, .EXTU7:focus, .UuUQYe:focus { outline: none; background-color: rgb(241, 243, 244); }

.UuUQYe { border-radius: 18px; flex: 0 0 auto; font-size: 0px; background-color: transparent; border: none; box-sizing: content-box; height: 18px; }

.rv4TOb { width: 18px; height: 18px; opacity: 0.55; }

.EXTU7 .rv4TOb { vertical-align: top; position: relative; top: -1px; }

.UuUQYe:hover > .rv4TOb, .UuUQYe:focus > .rv4TOb, .EXTU7:hover .rv4TOb, .EXTU7:focus .rv4TOb { opacity: 0.9; }

.n8vK9c { padding-right: 4px; }

.qGdXAc { font-family: "Google Sans", sans-serif; font-size: 13px; font-weight: 500; color: rgb(95, 99, 104); height: 18px; white-space: nowrap; }

.Kjhbcb { vertical-align: top; }

.qGdXAc:hover, .qGdXAc:focus { color: rgb(32, 33, 36); }

.MwUX8 { align-items: center; background-color: rgb(249, 249, 249); border: 0.0625em solid rgb(186, 186, 186); border-radius: 0.2em; bottom: 0.1em; box-sizing: border-box; display: inline-flex; height: 1.1em; justify-content: center; margin-left: 0.3em; position: relative; width: 1.8em; }

.DQD9Vb { color: rgb(186, 186, 186); font-size: 0.6em; font-weight: bold; }

.wvGCSb.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { background-color: rgb(11, 87, 208); }

.wvGCSb.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.HB1eCd-UMrnmb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { border-color: rgb(11, 87, 208); }

.wvGCSb-efwuC { background-color: rgb(245, 245, 245); cursor: pointer; direction: ltr; position: relative; width: 240px; border: none; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px; border-radius: 2px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC { background-color: rgb(255, 255, 255); border: 1px solid rgba(60, 64, 67, 0.15); box-shadow: none; width: 282px; }

.HB1eCd-UMrnmb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC { min-width: 282px; width: calc(100% - 50px); max-width: calc(50ch + 24px); }

.HB1eCd-UMrnmb .wvGCSb-efwuC:hover { border-color: transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover { border-color: transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC-k4Qmrd, .HB1eCd-UMrnmb .wvGCSb-efwuC { border-radius: 8px; }

.wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC { cursor: default; }

.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-UMrnmb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover, .HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover { background-color: transparent; cursor: pointer; border: none; box-shadow: none; }

.wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb-efwuC-Nk0Zid, .wvGCSb-efwuC-Nk0Zid .HB1eCd-Bz112c { min-height: 24px; min-width: 24px; max-width: 24px; }

.HB1eCd-UMrnmb .wvGCSb-Nk0Zid-nUpftc.wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .wvGCSb-Nk0Zid-nUpftc.wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:not(.wvGCSb-pnL5fc-auswjd):hover .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_dark.svg"); }

.wvGCSb-efwuC:focus, .wvGCSb-efwuC:active { outline: 0px; }

.wvGCSb-efwuC-k4Qmrd { max-height: inherit; overflow: hidden auto; }

.wvGCSb-efwuC-bN97Pc { overflow: hidden auto; }

.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { border: none; display: none; padding: 8px; }

.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc.wvGCSb-UbLY0d-YPqjbf-BeDmAc { padding-top: 0px; }

.wvGCSb-efwuC .wvGCSb-UbLY0d-YPqjbf-BeDmAc { background: rgb(255, 255, 255); }

.wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { display: block; }

.wvGCSb-RDNXzf-P7Vtfd .wvGCSb-efwuC-k4Qmrd { background: rgb(237, 242, 250); }

.wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { display: block; height: 26px; }

.wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-c6xFrd { text-align: left; }

.wvGCSb-UbLY0d-YPqjbf-BeDmAc { padding-top: 0px; border-top: none !important; }

.wvGCSb-efwuC .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .wvGCSb-efwuC .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .wvGCSb-efwuC .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .wvGCSb-efwuC .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(119, 119, 119); font-size: 12px; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin-top: 8px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; letter-spacing: 0.3px; line-height: 16px; }

.wvGCSb-neVct-uNfmef .wvGCSb-efwuC { position: absolute; user-select: text; z-index: 500; }

.wvGCSb-neVct-uNfmef .wvGCSb-CTWaPd-ZiwkRe.wvGCSb-efwuC { z-index: 502; }

.wvGCSb-neVct-uNfmef .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC { z-index: 501; }

.wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC { box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; }

.wvGCSb-efwuC .wvGCSb-YPqjbf-aIWppb { margin-right: 10px; }

.HB1eCd-UMrnmb .wvGCSb-neVct-BvBYQ .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb.wvGCSb-JYA2rd-dHwMxe { background-color: rgb(0, 0, 0); }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-Bz112c-qE2ISc { margin-top: 1px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Bz112c-qE2ISc { margin-top: 4px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC:hover { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb-eKrold-VkLyEc, .wvGCSb-eKrold-DyVDA { color: rgb(17, 85, 204); font-size: 11px; margin: 0px 2px; }

.wvGCSb-eKrold-VkLyEc:hover, .wvGCSb-eKrold-DyVDA:hover { text-decoration: underline; cursor: pointer; }

.wvGCSb-YPqjbf-IbE0S { margin: 0px; }

.wvGCSb-YPqjbf-aIWppb { margin: 8px 7px 0px 0px; }

.wvGCSb-H9tDt-xtcdFb-JIbuQc-fmcmS-sM5MNb { padding: 8px 0px 0px; position: relative; }

.wvGCSb-eKrold-giiMnc-GMvhG-fmcmS { overflow-wrap: break-word; margin: 8px -8px 0px; padding: 8px 8px 4px; border-color: rgb(229, 229, 229); border-top-style: solid; border-top-width: 1px; color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; line-height: 16px; }

.wvGCSb-Vq7Udc .wvGCSb-lCdvJf-fj0AZd { background-color: rgba(140, 196, 116, 0.5); }

.wvGCSb-Vq7Udc .wvGCSb-gk6SMd-lCdvJf-fj0AZd { background-color: rgb(140, 196, 116); }

.wvGCSb-Vq7Udc:focus { outline: none; }

.wvGCSb-Vq7Udc, .wvGCSb-BxnCYe { border-top: none; border-right: none; border-left: none; border-image: initial; border-bottom: 1px solid rgb(229, 229, 229); padding: 3px 8px 5px; zoom: 1; background: rgb(245, 245, 245); position: static; }

.wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 6px; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc { background-color: rgb(255, 255, 255); border-bottom: none; border-top: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb .wvGCSb-BxnCYe { background-color: rgb(255, 255, 255); border-bottom: none; }

.HB1eCd-UMrnmb .wvGCSb-efwuC-YPqjbf-BeDmAc { background-color: rgb(255, 255, 255); border-bottom: none; border-top: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb .wvGCSb-BxnCYe { border-top: none; color: rgb(26, 115, 232); letter-spacing: 0.2px; margin: 0px 8px; padding: 0px; position: relative; text-align: center; align-items: center; display: flex; justify-content: center; }

.HB1eCd-UMrnmb .wvGCSb-BxnCYe:not([style*="display: none"]) + .wvGCSb-Vq7Udc:not([style*="display: none"]), .HB1eCd-UMrnmb .wvGCSb-BxnCYe:not([style*="display: none"]) ~ .wvGCSb-Vq7Udc[style*="display: none"] + .wvGCSb-Vq7Udc:not([style*="display: none"]) { border-top: none; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-Vq7Udc { padding: 8px 0px; margin: 0px 12px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { border-bottom: none; padding: 12px 12px 8px; margin: 0px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 12px; }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-LgbsSe-oKdM2c { padding-top: 8px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.wvGCSb-efwuC .wvGCSb-efwuC-bN97Pc > .wvGCSb-Vq7Udc:last-of-type, .wvGCSb-efwuC .wvGCSb-pnL5fc-C58Yv:only-child .wvGCSb-Vq7Udc { padding-bottom: 12px; }

.wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { padding: 8px; border-bottom: 1px solid rgb(221, 221, 221); background: rgb(255, 255, 255); min-height: 36px; }

.wvGCSb-pnL5fc-IIEkAe .wvGCSb-Vq7Udc, .wvGCSb-pnL5fc-IIEkAe .wvGCSb-BxnCYe, .wvGCSb-efwuC.wvGCSb-pnL5fc-IIEkAe .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc, .HB1eCd-UMrnmb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-efwuC { background: rgb(238, 238, 238); }

.wvGCSb-efwuC .wvGCSb-efwuC-yqoORe .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { border: none; }

.wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-YLEF4c { display: block; left: 0px !important; }

.wvGCSb-Vq7Udc.wvGCSb-eKrold-r08add { border-top: none !important; }

.wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { margin: 2px 0px 0px; color: rgb(51, 51, 51); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; font-weight: 500; height: 18px; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { color: rgb(60, 64, 67); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; margin-top: 0px; }

.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od, .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM .wvGCSb-Vq7Udc-FDWhSe { line-height: 1.4; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { line-height: 20px; }

.wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { overflow-wrap: break-word; color: rgb(51, 51, 51); padding: 0px; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { color: rgb(0, 0, 0); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; letter-spacing: 0.2px; line-height: 20px; }

.wvGCSb-Vq7Udc .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy { padding: 3px 21px 3px 5px; }

.wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc { background-color: rgb(241, 243, 244); border-radius: 6px; }

.wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background: white; border-radius: 50%; bottom: -3px; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; display: flex; justify-content: center; padding: 0px; position: absolute; right: -14px; width: 32px; z-index: 10; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM a { color: rgb(26, 115, 232); }

.wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { margin: 0px; color: rgb(119, 119, 119); font-size: 11px; }

.HB1eCd-UMrnmb .QpLw9-qnnXGd-lI7fHe .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { align-items: center; display: inline-flex; flex-direction: row; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; letter-spacing: 0.3px; }

.HB1eCd-UMrnmb .wvGCSb-pnL5fc-MGbz6c .wvGCSb-RmniWd-mQXP { flex: 0 0 auto; align-items: center; background-color: rgb(26, 115, 232); border-radius: 9px; color: white; height: 16px; justify-content: center; margin: auto 0px; overflow: hidden; transform-origin: left center; transition: transform 0.2s ease-out 0s, color 0.1s ease-in 0s, border-radius 0.2s ease 0s; }

.HB1eCd-UMrnmb .wvGCSb-pnL5fc-MGbz6c:not(:hover) .wvGCSb-RmniWd-mQXP { border-radius: 50%; color: white; width: 6px; transform: scale(0.375); }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc span + .wvGCSb-RmniWd-mQXP { margin-left: 4px; }

.wvGCSb-RmniWd-mQXP { font-weight: 600; display: inline-block; font-size: 0.75rem; font-family: Roboto, sans-serif; padding: 0px 5px; }

.HB1eCd-UMrnmb .wvGCSb-pnL5fc-MGbz6c:not(:hover) .wvGCSb-RmniWd-Ne3sFf { color: transparent; }

.wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { min-width: 28px; width: 28px; }

.wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd { height: 28px; margin: 0px; position: relative; top: auto; display: inline-block; vertical-align: middle; }

.wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { height: 28px; margin: 0px; position: relative; top: auto; right: auto; display: inline-block; vertical-align: middle; }

.wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { padding: 0px; }

.wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd { right: -1px; }

.wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd div, .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd div { margin: 1px auto auto; }

.wvGCSb-no16zc-ldDtVd { border-radius: 3px 0px 0px 3px; }

.wvGCSb-ERydpb-ldDtVd { border-radius: 0px 3px 3px 0px; }

.wvGCSb.HB1eCd-UMrnmb .wvGCSb-no16zc-ldDtVd path, .wvGCSb.HB1eCd-UMrnmb .wvGCSb-ERydpb-ldDtVd path { fill: rgb(0, 0, 0); }

.wvGCSb.HB1eCd-UMrnmb .wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me path, .wvGCSb.HB1eCd-UMrnmb .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me path { fill: rgb(60, 64, 67); }

.wvGCSb.HB1eCd-UMrnmb .wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me, .wvGCSb.HB1eCd-UMrnmb .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me { background-color: white; opacity: 0.38; }

.wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me, .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me { background-color: rgb(249, 249, 249); }

.wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC .wvGCSb-eKrold-bMcfAe, .wvGCSb-pnL5fc-auswjd.wvGCSb-BxnCYe .wvGCSb-eKrold-bMcfAe { display: block; }

.wvGCSb-BxnCYe-qAWA2 { overflow-wrap: break-word; color: rgb(17, 85, 204); }

.wvGCSb-BxnCYe-qAWA2:hover, .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2 { text-decoration: underline; }

.wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:hover { text-decoration: underline; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2 { position: relative; width: 100%; }

.wvGCSb-efwuC .wvGCSb-BxnCYe-RWgCYc { border-top: 1px solid rgb(218, 220, 224); height: 50%; position: absolute; top: 50%; width: 100%; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd { background-color: rgb(255, 255, 255); display: inline-block; margin: 0px 20px; padding: 0px 8px; position: relative; overflow-wrap: break-word; word-break: break-word; }

.wvGCSb-rM9Gsd-eKrold { position: relative; margin: 6px 0px; padding: 0px; }

.HB1eCd-UMrnmb .wvGCSb-rM9Gsd-eKrold { margin-bottom: 0px; }

.wvGCSb-rM9Gsd-eKrold.wvGCSb-rM9Gsd-eKrold-xFQqWe { margin: 0px; }

.wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold { height: 78px; overflow: hidden; }

.wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 81px; overflow: hidden; }

.wvGCSb-ti6hGc-z5C9Gb, .wvGCSb-ti6hGc-OCFbXc { color: rgb(17, 85, 204); display: none; opacity: 1; width: 100%; outline: none; }

.wvGCSb-ti6hGc-z5C9Gb:focus, .wvGCSb-ti6hGc-OCFbXc:focus { text-decoration: underline; }

.wvGCSb-ti6hGc-z5C9Gb { bottom: 0px; padding-top: 16px; position: absolute; right: 0px; }

.wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { cursor: pointer; font-size: 11px; }

.wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc { background: rgb(245, 245, 245); padding: 2px 0px; }

.wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { padding: 7px 0px 2px; }

.wvGCSb-efwuC .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-OCFbXc { background: rgb(255, 255, 255); }

.wvGCSb-ti6hGc-z5C9Gb:hover, .wvGCSb-ti6hGc-OCFbXc:hover { text-decoration: underline; }

.wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.wvGCSb-efwuC .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-UMrnmb .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb-qAWA2-eKrold > .wvGCSb-eKrold-TJEFFc > .wvGCSb-ti6hGc-z5C9Gb { display: block; }

.wvGCSb-qAWA2-eKrold > .wvGCSb-eKrold-TJEFFc { height: 100%; }

.wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc > .wvGCSb-ti6hGc-z5C9Gb { display: block; }

.wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 100%; overflow: hidden; }

.wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc { background: rgb(245, 245, 245); }

.wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-OCFbXc { background: rgb(255, 255, 255); }

.wvGCSb-Vq7Udc-tJHJj { margin: 6px 0px; height: 38px; white-space: nowrap; display: flex; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-tJHJj { margin-top: 0px; }

.wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-tJHJj { margin: 0px 0px 8px; }

.wvGCSb-efwuC-yqoORe .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-tJHJj { margin: 0px; }

.wvGCSb-Vq7Udc-UwkkNe { white-space: nowrap; }

.wvGCSb-efwuC:hover .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd, .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd, .wvGCSb-efwuC.wvGCSb-CTWaPd-ZiwkRe .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd { border: 1px solid rgba(255, 255, 255, 0.7); }

.wvGCSb-W3vEtb-n0tgWb .VIpgJd-xl07Ob { z-index: 600; }

.wvGCSb-Vq7Udc-UwkkNe:hover .wvGCSb-ERydpb-ldDtVd, .wvGCSb-Vq7Udc-UwkkNe:hover .wvGCSb-eKrold-WlKKfd-LgbsSe { border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.wvGCSb-Vq7Udc-UwkkNe > .wvGCSb-ERydpb-ldDtVd:hover, .wvGCSb-Vq7Udc-UwkkNe > .wvGCSb-eKrold-WlKKfd-LgbsSe:hover { border-top-right-radius: 2px; border-bottom-right-radius: 2px; }

.wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-UwkkNe { padding: 4px 0px 4px 4px; }

.wvGCSb-no16zc-ldDtVd { margin-right: -1px; }

.wvGCSb-Vq7Udc-fXZhbb { padding-left: 10px; overflow: hidden; white-space: nowrap; text-overflow: ellipsis; -webkit-box-flex: 1; flex-grow: 1; }

.QpLw9-qnnXGd-lI7fHe .wvGCSb-Vq7Udc-fXZhbb span { overflow: hidden; text-overflow: ellipsis; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-fXZhbb { display: flex; align-items: start; flex-direction: column; justify-content: center; }

.wvGCSb-Vq7Udc-fXZhbb > * { overflow: hidden; text-overflow: ellipsis; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-fXZhbb > * { align-self: stretch; }

.wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { max-width: 32px; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { height: 38px; margin-top: 2px; max-width: 36px; width: 36px; }

.wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { position: relative; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { margin-left: 2px; margin-top: 2px; }

.wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd { display: inline-block; margin: 0px; opacity: 0.2; position: relative; padding: 0px 4px; min-width: 50px; height: 28px; vertical-align: top; }

.HB1eCd-UMrnmb .wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: white; color: rgb(26, 115, 232); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb .wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd:hover { background: rgb(248, 251, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb .wvGCSb-eKrold-WlKKfd-LgbsSe { border-radius: 3px 0px 0px 3px; display: inline-block; margin: 1px auto auto; padding: 0px; position: relative; top: auto; right: auto; vertical-align: middle; width: 28px; height: 28px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC:hover .wvGCSb-eKrold-WlKKfd-LgbsSe, .HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-WlKKfd-LgbsSe { opacity: 1; }

.wvGCSb-Vq7Udc .wvGCSb-eKrold-DyVDA { margin-left: 0px; }

.wvGCSb-Vq7Udc-FDWhSe { overflow-wrap: break-word; color: rgb(119, 119, 119); margin: 8px -8px 0px; padding: 8px 8px 4px; border-color: rgb(229, 229, 229); border-top-style: solid; border-top-width: 1px; font-size: 11px; font-style: italic; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc-FDWhSe { color: rgb(128, 134, 139); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; }

.wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS { color: rgb(112, 112, 112); font-style: italic; overflow-wrap: break-word; }

.HB1eCd-UMrnmb .wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS { color: rgb(128, 134, 139); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; letter-spacing: 0.2px; line-height: 20px; }

.wvGCSb-JIbuQc-fmcmS-cGMI2b-sM5MNb { padding: 8px 0px 3px; position: relative; }

.wvGCSb-efwuC .wvGCSb-Vq7Udc:last-of-type .wvGCSb-JIbuQc-fmcmS-cGMI2b-sM5MNb { padding: 8px 0px 0px; }

.wvGCSb-eKrold-GyPgRd-sM5MNb { display: flex; flex-wrap: wrap; padding-top: 5px; }

.wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border: 1px solid rgba(60, 64, 67, 0.15); border-radius: 15px; margin: 1.5px; }

.wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-image: radial-gradient(ghostwhite, lavender); cursor: inherit; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { padding: 16px 16px 8px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-pnL5fc-C58Yv :only-child.wvGCSb-Vq7Udc { padding-bottom: 12px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC { background: transparent; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(243, 246, 252); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { border: none; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-k4Qmrd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { border-radius: 12px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od:focus, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-YPqjbf-BeDmAc.wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od:focus { background: rgb(255, 255, 255); border: 1px solid rgb(199, 199, 199); border-radius: 18px; color: rgb(31, 31, 31); font-family: "Google Sans", Roboto, sans-serif; padding: 8px 7px 8px 16px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { border-color: rgb(199, 199, 199); margin: 0px 16px; }

.wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-Vq7Udc, .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { border-color: rgb(199, 199, 199); margin: 0px; }

.wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-Vq7Udc { padding-left: 16px; padding-right: 16px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM a { color: rgb(11, 87, 208); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(231, 237, 248); box-shadow: none; }

.wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC:hover { background: transparent; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd:hover .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd:hover .wvGCSb-efwuC-YPqjbf-BeDmAc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(255, 255, 255); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-UwkkNe { opacity: 0; transition: opacity 250ms cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-WlKKfd-LgbsSe, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { border: none; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-no16zc-ldDtVd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ERydpb-ldDtVd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc-UwkkNe, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-Vq7Udc-UwkkNe { opacity: 1; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { color: rgb(31, 31, 31); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-F6aDIf .wvGCSb-dhWRR-biJjHb, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-JIbuQc-fmcmS { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; font-size: 12px; font-style: normal; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-H9tDt-xtcdFb-JIbuQc-fmcmS-sM5MNb { padding-bottom: 2px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd div, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd div { margin-top: 2px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 0px 0px 16px; }

.wvGCSb-RDNXzf-P7Vtfd .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 0px 16px 16px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe { margin: 0px 16px; background: none; color: rgb(68, 71, 70); font: 500 14px / 20px "Google Sans", Roboto, sans-serif; -webkit-font-smoothing: antialiased; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe-qAWA2 { background: none; color: rgb(68, 71, 70); font: 500 14px / 20px "Google Sans", Roboto, sans-serif; -webkit-font-smoothing: antialiased; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd { border-radius: 100px; margin: 0px 8px; padding: 2px 8px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(237, 242, 250); display: inline-block; position: relative; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(243, 246, 252); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd { color: rgb(11, 87, 208); text-decoration: none; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(231, 237, 248); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:hover { background-color: rgba(11, 87, 208, 0.08); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:focus, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:active { background-color: rgba(11, 87, 208, 0.12); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc { background-color: rgba(68, 71, 70, 0.08); border-radius: 8px; outline: transparent solid 1px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { box-shadow: rgba(0, 0, 0, 0.3) 0px 2px 3px, rgba(0, 0, 0, 0.15) 0px 6px 10px 4px; padding: 0px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border-color: rgb(199, 199, 199); margin: 2px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-XpnDCe { border-color: transparent; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 2px 6px 2px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-color: rgb(225, 227, 225); background-image: none; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(237, 242, 250); font-family: "Google Sans", Roboto, sans-serif; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(243, 246, 252); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(231, 237, 248); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-pnL5fc-auswjd.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { max-width: 34px; width: 34px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { margin: 0px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-UwkkNe { padding: 0px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold { height: 81px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 87px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-RmniWd-mQXP.wvGCSb-RmniWd-mQXP { background-color: rgb(11, 87, 208); font: 500 11px / 16px "Google Sans", Roboto, sans-serif; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-ti6hGc-OCFbXc { color: rgb(11, 87, 208); text-decoration: none; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM span, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-qJTHM .wvGCSb-eKrold-qJTHM span { color: rgb(68, 71, 70) !important; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-XpnDCe { padding: 0px; }

@media screen and (forced-colors: active) {
  .wvGCSb-Vq7Udc .wvGCSb-lCdvJf-fj0AZd, .wvGCSb-efwuC .wvGCSb-gk6SMd-lCdvJf-fj0AZd { background-color: highlight; color: highlighttext; }
  .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc, .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { outline: highlight solid 1px; }
}

.wvGCSb-itKi9e-Btuy5e-haAclf { width: fit-content; }

.wvGCSb-itKi9e-Btuy5e { cursor: pointer; display: flex; height: 18px; margin: 4px 0px 8px; outline: transparent solid 1px; }

.wvGCSb-itKi9e-Btuy5e.HB1eCd-Guievd-WqyaDf { border: 1px solid transparent; }

.wvGCSb-itKi9e-Btuy5e .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

docs-blue-tint-icon-cleanup .wvGCSb-itKi9e-Btuy5e .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb-itKi9e-Btuy5e-fmcmS { color: rgb(26, 115, 232); font: 500 14px "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 0px 8px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e { align-items: center; border-radius: 12px; height: 24px; padding: 2px 8px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:hover { background: rgba(11, 87, 208, 0.08); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:focus, .HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:active { background: rgba(11, 87, 208, 0.12); }

.wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf .wvGCSb-gkA7Yd-Wz3zdc-T3yXSc-cHYyed { line-height: 20px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-style: normal; font-size: 14px; }

.wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(241, 243, 244); display: flex; flex-direction: row; align-items: center; padding: 10px 16px; border-top-left-radius: 8px; border-top-right-radius: 9px; margin: -1px; }

.wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc-JIbuQc-haAclf { display: flex; flex-direction: row; position: relative; padding-bottom: 15px; }

.wvGCSb-gkA7Yd-Wz3zdc-FDWhSe { color: rgb(128, 134, 139); font-size: 11px; font-style: italic; text-align: left; white-space: pre-wrap; }

.gkA7Yd-Wz3zdc-lI7fHe-nUpftc-tJHJj-clz4Ic { padding: 0px 5px; }

:not(docos-docoview-resolved) .wvGCSb-dhWRR:hover .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(254, 239, 195); }

:not(docos-docoview-resolved) .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(253, 214, 99); }

.wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf, .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(218, 220, 224); }

.wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc, .wvGCSb-pnL5fc-IIEkAe.wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc { background-color: rgb(241, 243, 244); }

.wvGCSb-gkA7Yd-Wz3zdc-MZArnb { position: absolute; right: 0px; top: 0px; }

.wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { display: none; }

.wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { margin: 0px 8px 0px 0px; width: 28px; height: 28px; vertical-align: middle; }

.wvGCSb-W3vEtb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { min-width: 14px; }

.wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc-j4LONd-cnfHN { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 18px; letter-spacing: 0.25px; line-height: 20px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-MZArnb { display: flex; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { align-items: center; display: flex; justify-content: center; background: none; border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb-F9IAbd-xtcdFb { display: flex; justify-content: space-between; text-align: center; margin-right: 6px; }

.wvGCSb.HB1eCd-UMrnmb .wvGCSb-F9IAbd-xtcdFb-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe { align-items: center; display: flex; height: auto; justify-content: center; padding: 3px 12px; white-space: normal; width: 100%; }

.wvGCSb-F9IAbd-xtcdFb .wvGCSb-F9IAbd-xtcdFb-LgbsSe:last-child { margin-right: 0px; }

.wvGCSb-F9IAbd-xtcdFb-LgbsSe-cHYyed { display: inline; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .wvGCSb-F9IAbd-xtcdFb .wvGCSb-F9IAbd-xtcdFb-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe { border-radius: 18px; height: auto; min-height: 36px; padding: 3px 12px; }

.wvGCSb-YPqjbf { position: relative; outline: none; zoom: 1; }

.wvGCSb-YPqjbf.wvGCSb-YPqjbf-mOyJmb { display: block !important; }

.wvGCSb-YPqjbf-lvBGLe { cursor: text; text-align: start; overflow-wrap: break-word; }

.wvGCSb-YPqjbf-lvBGLe:empty::before { color: rgb(128, 134, 139); content: attr(placeholder); display: block; pointer-events: none; }

@media screen and (forced-colors: active) {
  .wvGCSb-YPqjbf-lvBGLe:empty::before { color: graytext; }
}

.wvGCSb-YPqjbf-lvBGLe p { margin: 0px; }

.wvGCSb-YPqjbf-B7I4Od { box-sizing: border-box; color: rgb(153, 153, 153); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; margin: 0px; overflow: hidden; padding: 4px; resize: none; width: 100%; border: 1px solid rgb(200, 200, 200); outline-width: 0px !important; }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-B7I4Od { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(60, 64, 67); font-size: 14px; line-height: 20px; min-height: 36px; padding: 8px; }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-B7I4Od:focus { border: 2px solid rgb(26, 115, 232); box-shadow: none; padding: 7px; }

.wvGCSb-YPqjbf-B7I4Od:disabled { background-color: rgb(238, 238, 238) !important; }

:first-child + html .wvGCSb-YPqjbf-B7I4Od { width: 95%; }

.wvGCSb-YPqjbf-c6xFrd { display: none; zoom: 1; }

.wvGCSb-YPqjbf-c6xFrd-aIWppb { font-weight: 500; }

.wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { color: rgb(0, 0, 0); }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { color: rgb(60, 64, 67); }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { background-color: rgb(255, 255, 255); }

.wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-c6xFrd { display: block; }

.wvGCSb-YPqjbf-IIyL0-wcotoc-fmcmS { color: rgb(97, 97, 97); font-style: italic; padding: 5px 0px 3px; overflow-wrap: break-word; }

.wvGCSb-YPqjbf-lQVAed-b0t70b { padding: 6px 8px 4px; background-color: rgb(245, 245, 245); border-style: solid; border-width: 0px 1px 1px; border-color: rgb(200, 200, 200); margin-bottom: 8px; cursor: pointer; }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-lQVAed-b0t70b { padding: 6px 8px 11px 0px; background-color: rgb(255, 255, 255); border-width: 1px; border-style: solid; border-color: transparent transparent rgb(218, 220, 224); border-image: initial; margin-bottom: 18px; cursor: pointer; }

.wvGCSb-YPqjbf-lQVAed-Q4BLdf { margin: 2px 10px 0px 0px; float: left; width: 11px; }

.wvGCSb-efwuC .wvGCSb-YPqjbf-JYA2rd-fmcmS { margin-top: 1px; }

.wvGCSb-YPqjbf-JYA2rd-fmcmS { text-align: left; white-space: nowrap; overflow: hidden; text-overflow: ellipsis; font-size: 13px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(112, 112, 112); font-weight: normal; display: inline-block; width: calc(100% - 51px); }

.wvGCSb-YPqjbf-JYA2rd-fmcmS.wvGCSb-YPqjbf-JYA2rd-fmcmS-di8rgd-Q8Kwad { width: calc(100% - 23px); }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-JYA2rd-fmcmS { margin-top: 6px; margin-left: 8px; white-space: nowrap; overflow: hidden; text-overflow: ellipsis; font-size: 14px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(60, 64, 67); font-weight: normal; display: inline-block; width: calc(100% - 57px); }

.HB1eCd-UMrnmb .wvGCSb-YPqjbf-JYA2rd-fmcmS.wvGCSb-YPqjbf-JYA2rd-fmcmS-di8rgd-Q8Kwad { width: calc(100% - 29px); }

.wvGCSb-dhWRR .wvGCSb-YPqjbf-JYA2rd-O1htCb { margin-top: 0px; }

.wvGCSb-JYA2rd-O1htCb-AHmuwe { border-radius: 2px; border: 1px solid rgb(77, 144, 254) !important; }

.wvGCSb-YPqjbf-JYA2rd-O1htCb { border: none; background: none; box-shadow: none; cursor: pointer; float: right; width: 24px; height: 15px; margin: 2px; }

.HB1eCd-UMrnmb .wvGCSb-efwuC .wvGCSb-YPqjbf-JYA2rd-O1htCb { margin-top: 6px; }

.wvGCSb-YPqjbf-JYA2rd-O1htCb .VIpgJd-xl07Ob-LgbsSe-cHYyed { padding: 0px; }

.wvGCSb-YPqjbf-JYA2rd-O1htCb .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { margin: 0px; }

.wvGCSb-JYA2rd-O1htCb-ibnC6b { padding: 0px; border-width: 0px; }

.wvGCSb-JYA2rd-O1htCb-ibnC6b.VIpgJd-j7LFlb-sn54Q { background-color: rgb(242, 242, 242); }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.wvGCSb-JYA2rd-O1htCb-xl07Ob { padding: 4px 0px; max-height: 222px; overflow-y: auto; box-sizing: border-box; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob { padding: 8px 0px; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob .wvGCSb-JYA2rd-O1htCb-ibnC6b, .VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob .wvGCSb-JYA2rd-O1htCb-ibnC6b.VIpgJd-xl07Ob-ibnC6b-sn54Q { border: none; padding: 0px; }

.wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-j4gsHd { width: 24px; background: url("//ssl.gstatic.com/images/icons/material/system/2x/arrow_drop_down_black_24dp.png") center center / 24px no-repeat; opacity: 0.54; box-sizing: border-box; }

.wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-j4gsHd:hover { opacity: 0.87; }

.wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-style: none; padding: 0px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf-lvBGLe:empty::before { color: rgb(68, 71, 70); }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf-lQVAed-b0t70b { background-color: inherit; }

.tk3N6e-MPu53c { border-radius: 1px; background-color: rgba(255, 255, 255, 0.05); border: 1px solid rgba(155, 155, 155, 0.57); font-size: 1px; height: 11px; margin: 0px 4px 0px 1px; outline: 0px; vertical-align: text-bottom; width: 11px; }

.tk3N6e-MPu53c-uE9yNd, .tk3N6e-MPu53c-barxie { background-color: rgba(255, 255, 255, 0.65); }

.tk3N6e-MPu53c-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px inset; border: 1px solid rgb(178, 178, 178); }

.tk3N6e-MPu53c-auswjd { background-color: rgb(235, 235, 235); }

.tk3N6e-MPu53c-XpnDCe { border: 1px solid rgb(77, 144, 254); }

.tk3N6e-MPu53c-kyhDef.tk3N6e-MPu53c-XpnDCe { border: 1px solid rgba(155, 155, 155, 0.57); }

.tk3N6e-MPu53c-OWB6Me, .tk3N6e-MPu53c-kyhDef.tk3N6e-MPu53c-OWB6Me { background-color: rgb(255, 255, 255); border: 1px solid rgb(241, 241, 241); cursor: default; }

.tk3N6e-MPu53c-qE2ISc { height: 15px; outline: 0px; width: 15px; left: 0px; position: relative; top: -3px; }

.tk3N6e-MPu53c-uE9yNd .tk3N6e-MPu53c-qE2ISc { background: image-set(url("//ssl.gstatic.com/ui/v1/menu/checkmark-partial.png") 1x, url("//ssl.gstatic.com/ui/v1/menu/checkmark-partial_2x.png") 2x) -5px -3px no-repeat; }

.tk3N6e-MPu53c-barxie .tk3N6e-MPu53c-qE2ISc { background: image-set(url("//ssl.gstatic.com/ui/v1/menu/checkmark.png") 1x, url("//ssl.gstatic.com/ui/v1/menu/checkmark_2x.png") 2x) -5px -3px no-repeat; }

.Jiyx5 { list-style: none; margin: 0px; padding: 0px; }

.Jiyx5:focus { outline: none; }

.MsdWL { background: rgb(255, 255, 255); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.aqWPhc .MsdWL { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.MsdWL.nhiZfc { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; height: 48px; }

.MsdWL.nhiZfc .E8WqE { height: 24px; width: 24px; margin-right: 16px; }

.MsdWL.XdSAtd { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; height: 32px; }

.MsdWL.XdSAtd .E8WqE { height: 20px; width: 20px; margin-right: 12px; }

.MsdWL.HddOwd { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; height: 32px; }

.MsdWL.HddOwd .E8WqE { height: 20px; width: 20px; margin-right: 12px; }

.MsdWL:hover { background: rgba(10, 10, 10, 0.04); }

.aqWPhc .MsdWL:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.MsdWL.qs41qe { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; }

.aqWPhc .MsdWL.qs41qe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.25), rgba(232, 234, 237, 0.25)), rgb(32, 33, 36); }

.jcbibd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; max-width: 450px; padding-left: 12px; padding-right: 12px; }

.w8bLS { -webkit-box-flex: initial; flex: initial; }

.B92god { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.hMC4ff { -webkit-box-flex: initial; flex: initial; }

.E8WqE { margin-left: 0px; }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .E8WqE { filter: brightness(0) invert(1); }
}

.EKzqb { color: rgb(60, 64, 67); text-overflow: ellipsis; white-space: nowrap; }

.aqWPhc .EKzqb { color: rgb(232, 234, 237); }

.bylmg { color: rgb(95, 99, 104); margin-left: 48px; margin-right: 0px; white-space: nowrap; }

.aqWPhc .bylmg { color: rgb(218, 220, 224); }

.heO6Yc { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 4px; outline: transparent solid 1px; overflow: hidden; padding-bottom: 8px; padding-top: 8px; position: absolute; user-select: none; z-index: 999999; }

.heO6Yc .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.aqWPhc .heO6Yc { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.O5UuBc { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; color: rgb(26, 115, 232); -webkit-box-align: center; align-items: center; background: none; border-radius: 4px; border: none; outline: transparent solid 1px; display: flex; height: 36px; line-height: unset; padding: 0px 8px; user-select: none; }

.aqWPhc .O5UuBc { color: rgb(138, 180, 248); }

.O5UuBc:hover { background-color: rgba(26, 115, 232, 0.04); color: rgb(23, 78, 166); cursor: pointer; }

.aqWPhc .O5UuBc:hover { background-color: rgba(138, 180, 248, 0.04); color: rgb(210, 227, 252); }

.O5UuBc:focus { background-color: rgba(26, 115, 232, 0.12); color: rgb(23, 78, 166); cursor: pointer; outline-width: 3px; }

.aqWPhc .O5UuBc:focus { background-color: rgba(138, 180, 248, 0.12); color: rgb(210, 227, 252); }

.O5UuBc.RDPZE { color: rgba(60, 64, 67, 0.38); }

.aqWPhc .O5UuBc.RDPZE { color: rgba(232, 234, 237, 0.38); }

.O5UuBc.RDPZE:focus { background-color: rgba(60, 64, 67, 0.12); color: rgba(60, 64, 67, 0.38); }

.aqWPhc .O5UuBc.RDPZE:focus { background-color: rgba(232, 234, 237, 0.12); color: rgba(232, 234, 237, 0.38); }

.q5Gute { -webkit-box-align: center; align-items: center; background: rgba(32, 33, 36, 0.6); box-sizing: border-box; display: flex; height: 100%; -webkit-box-pack: center; justify-content: center; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 999999; }

.qnxR0c { background: rgb(255, 255, 255); }

.aqWPhc .qnxR0c { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.cySkyb { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 8px; max-width: 300px; outline: transparent solid 1px; overflow: hidden; }

.cySkyb .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.aqWPhc .cySkyb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.h6zUze { margin: 24px 24px 20px; }

.tAzG6 { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 8px; }

.g9hvRc { width: 8px; }

.xQiMxd { -webkit-box-align: center; align-items: center; background: rgba(32, 33, 36, 0.6); box-sizing: border-box; display: flex; height: 100%; -webkit-box-pack: center; justify-content: center; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 999999; }

.mSjfjb { background: rgb(255, 255, 255); }

.aqWPhc .mSjfjb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.tFDhVb { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 500; color: rgb(32, 33, 36); margin: 24px 24px 20px; }

.aqWPhc .tFDhVb { color: rgb(232, 234, 237); }

.EoolDb { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 8px; max-width: 300px; outline: transparent solid 1px; overflow: hidden; }

.EoolDb .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.aqWPhc .EoolDb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.Pmtn0b { margin: 24px 24px 20px; }

.X23yUb { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(60, 64, 67); margin-bottom: 24px; }

.aqWPhc .X23yUb { color: rgb(232, 234, 237); }

.ADqTKb { color: rgb(26, 115, 232); text-decoration: underline; white-space: nowrap; }

.aqWPhc .ADqTKb { color: rgb(138, 180, 248); }

.ADqTKb:visited { color: rgb(26, 115, 232); }

.aqWPhc .ADqTKb:visited { color: rgb(138, 180, 248); }

.tlQjad { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 8px; }

.mtq6kd { position: relative; }

.A6DTme { border-radius: 50%; outline: transparent solid 1px; overflow: hidden; }

.hIJ6Le { margin: auto; display: block; height: 100%; width: 100%; }

.vi1cfb { position: absolute; bottom: 0px; right: 0px; display: none; height: 30%; width: 30%; min-height: 30%; min-width: 30%; object-fit: cover; overflow: hidden; }

.vi1cfb.ZiwkRe { display: inline; }

.KKjvXb .vi1cfb { display: none; }

.PS6m6 { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; height: inherit; width: inherit; }

.aGbmDb { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 0%; overflow: hidden; height: inherit; -webkit-box-align: stretch; align-items: stretch; }

.AcwQxb { display: flex; -webkit-box-flex: 1; flex: 1 1 0%; overflow: hidden; }

.IW1j2d { margin: 1px; }

.Khf4w { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 auto; -webkit-box-align: center; place-items: center; transition: background 50ms ease-in-out 0s; }

.Khf4w.JpY6Fd { background-clip: padding-box; background-color: rgb(189, 193, 198); }

.ew7bve { display: none; }

.k8rr2e .ew7bve { display: block; fill: rgb(95, 99, 104); }

.aqWPhc .k8rr2e .ew7bve { fill: rgb(154, 160, 166); }

.ZlXryd { opacity: 1; display: block; transition: opacity 50ms ease-in-out 0s; }

.JpY6Fd .ZlXryd { opacity: 0; }

.k8rr2e .ZlXryd { display: none; }

.AGaBze { background: rgb(255, 255, 255); border-bottom: 1px solid rgb(218, 220, 224); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.aqWPhc .AGaBze { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.haq1x { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; padding: 12px; }

.rr5U0b { -webkit-box-flex: initial; flex: initial; }

.tJRcje { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.XsnHSd { align-content: flex-start; -webkit-box-align: start; align-items: flex-start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-flow: column nowrap; margin-left: 12px; margin-right: 0px; }

.RWXYif { -webkit-box-flex: initial; flex: initial; width: 100%; }

.awj5uc { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; color: rgb(32, 33, 36); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.aqWPhc .awj5uc { color: rgb(232, 234, 237); }

.J7kVrb { font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; color: rgb(60, 64, 67); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.aqWPhc .J7kVrb { color: rgb(154, 160, 166); }

.fasgab { position: relative; }

.vG6Gfe { height: inherit; position: relative; width: inherit; }

.L7D8v { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; }

.aAzAef { margin-bottom: 20px; font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(32, 33, 36); }

.aqWPhc .aAzAef { color: rgb(255, 255, 255); }

.TeNodb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; color: rgb(60, 64, 67); margin-bottom: 24px; }

.aqWPhc .TeNodb { color: rgb(232, 234, 237); }

.AZW99 { background: rgb(255, 255, 255); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; cursor: pointer; }

.aqWPhc .AZW99 { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.AZW99.nhiZfc { height: 64px; }

.AZW99.nhiZfc .rNlsc { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; }

.AZW99.nhiZfc .O7pQ4 { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; }

.AZW99.nhiZfc .bRdBfe { width: 24px; height: 24px; }

.AZW99.nhiZfc .DcfYrb { width: 25px; height: 25px; }

.AZW99.nhiZfc .kcuFCe { padding-left: 16px; padding-right: 16px; }

.AZW99.XdSAtd { height: 52px; }

.AZW99.XdSAtd .rNlsc { font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; line-height: 1.25rem; }

.AZW99.XdSAtd .O7pQ4 { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; line-height: 1rem; }

.AZW99.XdSAtd .bRdBfe { width: 19px; height: 19px; }

.AZW99.XdSAtd .DcfYrb { width: 20px; height: 20px; }

.AZW99.XdSAtd .kcuFCe { padding-left: 12px; padding-right: 12px; }

.AZW99.HddOwd { height: 44px; }

.AZW99.HddOwd .rNlsc { font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; line-height: 1.125; }

.AZW99.HddOwd .O7pQ4 { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; line-height: 0.875rem; }

.AZW99.HddOwd .bRdBfe { width: 17px; height: 17px; }

.AZW99.HddOwd .DcfYrb { width: 20px; height: 20px; }

.AZW99.HddOwd .kcuFCe { padding-left: 12px; padding-right: 12px; }

.AZW99.RDPZE { cursor: default; }

.AZW99.RDPZE .rNlsc, .AZW99.RDPZE .G1zVib { color: rgb(60, 64, 67); opacity: 0.38; }

.aqWPhc .AZW99.RDPZE .rNlsc, .aqWPhc .AZW99.RDPZE .G1zVib { color: rgb(232, 234, 237); }

.AZW99.RDPZE .p1rXue { opacity: 0.5; }

.AZW99.KKjvXb .s38Kwb { opacity: 1; transform: scale(1); }

.AZW99:hover { background: rgba(10, 10, 10, 0.04); }

.aqWPhc .AZW99:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.AZW99.qs41qe { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.aqWPhc .AZW99.qs41qe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.AZW99.FdSZEb { background-color: papayawhip; }

.kcuFCe { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; }

.r6EVzf { -webkit-box-flex: initial; flex: initial; }

.uy8S0e { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.arWWkb { display: inline-flex; -webkit-box-flex: initial; flex: initial; }

.CnoS1b { align-content: flex-start; -webkit-box-align: start; align-items: flex-start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-flow: column nowrap; margin-left: 12px; margin-right: 0px; }

.pX5gAc { -webkit-box-flex: initial; flex: initial; width: 100%; }

.rNlsc { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.PNwDub { color: rgb(60, 64, 67); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.aqWPhc .PNwDub { color: rgb(232, 234, 237); }

.dUj0G { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-align: center; align-items: center; }

.O7pQ4 { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.G1zVib { color: rgb(95, 99, 104); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.aqWPhc .G1zVib { color: rgb(154, 160, 166); }

.p1rXue { position: relative; }

.wRSMoe { height: inherit; width: inherit; position: relative; }

.s38Kwb { background-color: rgb(26, 115, 232); border-radius: 50%; height: 100%; left: 0px; opacity: 0; outline: transparent solid 1px; position: absolute; top: 0px; transform: scale(0); transition: transform 0.15s ease-out 0s, -webkit-transform 0.15s ease-out 0s; width: 100%; display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; }

.aqWPhc .s38Kwb { background-color: rgb(138, 180, 248); }

.GeKaSb { fill: rgb(255, 255, 255); display: inline-flex; }

.aqWPhc .GeKaSb { fill: rgb(32, 33, 36); }

@media (forced-colors: active) and (prefers-color-scheme: light) {
  .GeKaSb { filter: invert(1); }
}

.Hcawbb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; color: rgb(95, 99, 104); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; display: none; }

.DcfYrb { margin-left: 16px; margin-right: 4px; }

.DcfYrb[src=""] { display: none; }

.S3hTZb { background-color: rgb(241, 243, 244); color: rgb(32, 33, 36); display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-align: center; align-items: center; margin-left: 8px; border-radius: 4px; outline: transparent solid 1px; overflow: hidden; }

.S3hTZb.rNe0id { background-color: rgb(251, 188, 4); color: rgb(32, 33, 36); }

.nhiZfc .S3hTZb { height: 20px; min-width: 20px; }

.XdSAtd .S3hTZb, .HddOwd .S3hTZb { height: 16px; min-width: 16px; }

.nhiZfc .iHLOxc { width: 16px; height: 16px; margin-left: 2px; }

.XdSAtd .iHLOxc, .HddOwd .iHLOxc { width: 14px; height: 14px; margin-left: 1px; }

.R8dRld { max-width: 0px; overflow: hidden; transition: max-width 0.3s ease 0s; }

.S3hTZb:hover .R8dRld { max-width: 1000px; }

.xvZBXb { margin-left: 4px; margin-right: 4px; }

.nhiZfc .xvZBXb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; }

.XdSAtd .xvZBXb, .HddOwd .xvZBXb { font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; }

.KMIgo { -webkit-box-align: center; align-items: center; display: flex; }

.US5TTd { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(95, 99, 104); }

.aqWPhc .US5TTd { color: rgb(255, 255, 255); }

.l71Ouc { display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; background-color: rgb(241, 243, 244); border-radius: 50px; width: 32px; height: 32px; margin-left: 16px; margin-right: 4px; }

.aqWPhc .l71Ouc { background-color: rgba(241, 243, 244, 0.14); }

.LYstE { fill: rgb(95, 99, 104); }

.aqWPhc .LYstE { fill: rgb(232, 234, 237); }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .LYstE { filter: brightness(0) invert(1); }
}

.IYrrvc { background: none; border: none; border-radius: 50%; cursor: pointer; }

.IYrrvc:hover { background-color: rgb(218, 220, 224); }

.aqWPhc .IYrrvc:hover { background-color: rgb(95, 99, 104); }

.IYrrvc:active { background-color: rgb(189, 193, 198); }

.aqWPhc .IYrrvc:active { background-color: rgb(128, 134, 139); }

.IYrrvc.u3bW4e { background-color: rgb(218, 220, 224); outline: transparent solid 3px; }

.aqWPhc .IYrrvc.u3bW4e { background-color: rgb(95, 99, 104); }

.IYrrvc.nhiZfc { height: 40px; padding: 8px; width: 40px; }

.IYrrvc.nhiZfc .ssmXx { height: 24px; width: 24px; }

.IYrrvc.XdSAtd { height: 32px; padding: 6px; width: 32px; }

.IYrrvc.XdSAtd .ssmXx { height: 20px; width: 20px; }

.IYrrvc.HddOwd { height: 28px; padding: 5px; width: 28px; }

.IYrrvc.HddOwd .ssmXx { height: 18px; width: 18px; }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .IYrrvc .ssmXx { filter: brightness(0) invert(1); }
}

.L5nWEe { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; background-color: rgb(60, 64, 67); color: rgb(241, 243, 244); border-radius: 5px; box-sizing: border-box; line-height: 16px; min-width: 40px; max-width: 200px; min-height: 24px; max-height: 40vh; overflow: hidden; padding: 4px 8px; position: fixed; outline: transparent solid 1px; text-align: center; font-weight: bold; width: max-content; z-index: 9; }

.aqWPhc .L5nWEe { background-color: rgb(60, 64, 67); color: rgb(232, 234, 237); }

.hxyQfd { -webkit-box-align: center; align-items: center; border-radius: 50%; cursor: pointer; display: flex; transition: transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.hxyQfd:hover { background: rgba(10, 10, 10, 0.04); }

.aqWPhc .hxyQfd:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.hxyQfd:active { background: rgba(10, 10, 10, 0.12); }

.aqWPhc .hxyQfd:active { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.hxyQfd.TICPrf { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.aqWPhc .hxyQfd.TICPrf { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.hxyQfd.ReqAjb { transform: rotate(-180deg); }

.e63afb { fill: rgb(95, 99, 104); }

.aqWPhc .e63afb { fill: rgb(241, 243, 244); }

.EhtNt { -webkit-box-align: center; align-items: center; border-radius: 50%; cursor: pointer; display: flex; transition: transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.EhtNt:hover { background: rgba(10, 10, 10, 0.04); }

.aqWPhc .EhtNt:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.EhtNt:active { background: rgba(10, 10, 10, 0.12); }

.aqWPhc .EhtNt:active { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.EhtNt.TICPrf { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.aqWPhc .EhtNt.TICPrf { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.LGD9cb { fill: rgb(95, 99, 104); height: 16px; padding: 5px; width: 16px; }

.aqWPhc .LGD9cb { fill: rgb(241, 243, 244); }

.XhBoVe { background: rgb(255, 255, 255); }

.aqWPhc .XhBoVe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.a2oM9e { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; padding-left: 16px; padding-right: 16px; }

.TUsLr { color: rgb(95, 99, 104); font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.6875rem; letter-spacing: 0.0727273em; font-weight: 500; text-transform: uppercase; padding-bottom: 12px; padding-top: 12px; }

.aqWPhc .TUsLr { color: rgb(241, 243, 244); }

.xvJ2yc { flex-shrink: initial; flex-basis: initial; -webkit-box-flex: 1; flex-grow: 1; }

.xAiMkd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-pack: justify; justify-content: space-between; }

.F2iRTc { -webkit-box-flex: initial; flex: initial; }

.GZQpmf { -webkit-box-flex: initial; flex: initial; margin-left: 16px; margin-right: 4px; }

.RWYkoe { overflow: hidden; transform-origin: center top; transition: all 0.5s cubic-bezier(0.05, 0.7, 0.1, 1) 0s; }

.RWYkoe.qAWA2 { height: 0px; transform: scaleY(0); transition: all 0.2s cubic-bezier(0.3, 0, 0.8, 0.15) 0s; }

.FDlMAe { background: rgb(255, 255, 255); color: rgb(95, 99, 104); font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.6875rem; letter-spacing: 0.0727273em; font-weight: 500; text-transform: uppercase; padding-bottom: 12px; padding-left: 16px; padding-top: 12px; }

.aqWPhc .FDlMAe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); color: rgb(241, 243, 244); }

.pIQtMd { background: rgb(255, 255, 255); height: 100%; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; user-select: none; }

.aqWPhc .pIQtMd { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.pIQtMd.JpY6Fd .L5WGxc, .pIQtMd.JpY6Fd .zcyXfd { display: none; }

.pIQtMd.JpY6Fd .z7ZqLc { display: flex; -webkit-box-pack: center; justify-content: center; -webkit-box-align: center; align-items: center; height: 100%; }

.pIQtMd.JpY6Fd .z7ZqLc::before { -webkit-box-flex: 1; flex: 1 1 auto; }

.pIQtMd.JpY6Fd .z7ZqLc::after { -webkit-box-flex: 1; flex: 1 1 auto; }

.pIQtMd.Cn4kwe .L5WGxc, .pIQtMd.Cn4kwe .z7ZqLc { display: none; }

.pIQtMd.Cn4kwe .zcyXfd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: start; justify-content: flex-start; -webkit-box-align: center; align-items: center; height: 100%; overflow: auto; }

.L5WGxc { height: 100%; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; }

.z7ZqLc, .zcyXfd { display: none; }

.MFfTvd { display: inline-block; height: 40px; position: relative; width: 40px; direction: ltr; }

.FxUiNc { height: 0px; overflow: hidden; position: absolute; width: 0px; }

.QPPI1e { width: 100%; height: 100%; }

.MFfTvd.qs41qe .QPPI1e { animation: 1568ms linear 0s infinite normal none running circular-progress-container-rotate; }

.KLPWzf { height: 100%; opacity: 0; position: absolute; width: 100%; }

.Y6U90b { border-color: rgb(66, 133, 244); }

.l36Xze { border-color: rgb(234, 67, 53); }

.GybXwf { border-color: rgb(251, 188, 4); }

.v5iurb { border-color: rgb(52, 168, 83); }

.MFfTvd.qs41qe .KLPWzf.Y6U90b { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-blue-fade-in-out; }

.MFfTvd.qs41qe .KLPWzf.l36Xze { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-red-fade-in-out; }

.MFfTvd.qs41qe .KLPWzf.GybXwf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-yellow-fade-in-out; }

.MFfTvd.qs41qe .KLPWzf.v5iurb { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-green-fade-in-out; }

.OEwgzc { position: absolute; box-sizing: border-box; top: 0px; left: 45%; width: 10%; height: 100%; overflow: hidden; border-color: inherit; }

.OEwgzc .z58N3b { width: 1000%; left: -450%; }

.tEVydc { display: inline-block; position: relative; width: 50%; height: 100%; overflow: hidden; border-color: inherit; }

.tEVydc .z58N3b { width: 200%; }

.z58N3b { position: absolute; inset: 0px; box-sizing: border-box; height: 100%; border-width: 3px; border-style: solid; border-top-color: inherit; border-right-color: inherit; border-left-color: inherit; border-bottom-color: transparent; border-radius: 50%; animation: 0s ease 0s 1 normal none running none; }

.tEVydc.A9Yu7d .z58N3b { border-right-color: transparent; transform: rotate(129deg); }

.tEVydc.scD29d .z58N3b { left: -100%; border-left-color: transparent; transform: rotate(-129deg); }

.MFfTvd.qs41qe .tEVydc.A9Yu7d .z58N3b { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-left-spin; }

.MFfTvd.qs41qe .tEVydc.scD29d .z58N3b { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-right-spin; }

.MFfTvd.sf4e6b .QPPI1e { animation: 1568ms linear 0s infinite normal none running circular-progress-container-rotate, 400ms cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running circular-progress-fade-out; }

@-webkit-keyframes circular-progress-container-rotate { 
  100% { transform: rotate(360deg); }
}

@keyframes circular-progress-container-rotate { 
  100% { transform: rotate(360deg); }
}

@-webkit-keyframes circular-progress-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@keyframes circular-progress-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(1080deg); }
}

@-webkit-keyframes circular-progress-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@keyframes circular-progress-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@-webkit-keyframes circular-progress-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@keyframes circular-progress-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@-webkit-keyframes circular-progress-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@keyframes circular-progress-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@-webkit-keyframes circular-progress-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes circular-progress-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@-webkit-keyframes circular-progress-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@keyframes circular-progress-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@-webkit-keyframes circular-progress-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@keyframes circular-progress-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@-webkit-keyframes circular-progress-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes circular-progress-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

.wZ7wOe { border: none; outline: none; overflow: auto; }

.wZ7wOe::-webkit-scrollbar-thumb { background: rgb(221, 221, 221); border-width: 1px 4px; border-style: solid; border-color: white; border-radius: 8px; box-shadow: none; min-height: 40px; }

.wZ7wOe::-webkit-scrollbar-thumb:active { background: rgb(95, 99, 104); }

.wZ7wOe:hover::-webkit-scrollbar-thumb, .wZ7wOe::-webkit-scrollbar-thumb:hover { background: rgb(128, 134, 139); }

.HJOG0e { color: rgb(95, 99, 104); padding: 2em; text-align: center; -webkit-box-align: center; align-items: center; }

.aqWPhc .HJOG0e { color: rgb(154, 160, 166); }

.E633ec { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 500; }

.LPP4B { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; }

.YlzPUb { color: inherit; text-decoration: underline; white-space: nowrap; }

.OFaVze { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 4px; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; outline: transparent solid 2px; overflow: hidden; padding-bottom: 8px; padding-top: 8px; position: absolute; user-select: none; z-index: 999999; }

.OFaVze .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.aqWPhc .OFaVze { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { display: flex; align-items: center; height: 100%; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { background-size: contain; height: 24px; width: 24px; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { font-family: "Noto Color Emoji", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 20px; height: 32px; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-NnAfwf { align-items: center; display: flex; font-size: 14px; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c-haAclf { display: flex; flex-direction: row; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf > * { padding: 0px 3px; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-dIxMhd-Ca9lu.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { color: rgb(26, 115, 232); font-weight: 500; }

:not(.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-dIxMhd-Ca9lu).HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { color: rgb(95, 99, 104); font-weight: 400; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-PrY1nf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c-haAclf { font-size: 18px; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc { background-color: rgb(255, 255, 255); border-radius: 8px; box-shadow: rgb(189, 193, 198) 1px 0px 8px 1px; color: rgb(95, 99, 104); display: flex; font-size: 13px; font-weight: 400; line-height: 20px; margin-top: 7px; max-width: 258px; padding: 4px; text-align: center; width: auto; }

.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG, .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-color: rgb(255, 255, 255) transparent; left: -6px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { height: 32px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { align-items: center; display: flex; justify-content: center; width: 100%; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb.HB1eCd-HzV7m-LgbsSe { height: 24px; padding: 0px 5px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { height: 20px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { font-size: 16px; }

.HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf > * { padding: 0px 1px; }

.wvGCSb-PLt2Ue-haAclf { line-height: 140%; outline: none; }

.wvGCSb-PLt2Ue-bN97Pc { position: relative; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-PLt2Ue-bN97Pc { position: static; }

.wvGCSb-PLt2Ue-XHP5j { color: rgb(17, 85, 204); cursor: pointer; font-size: 12px; position: absolute; right: 0px; top: -3px; }

.wvGCSb-PLt2Ue-XHP5j:hover { text-decoration: underline; }

.wvGCSb-PrY1nf .wvGCSb-PLt2Ue-XHP5j { color: rgb(153, 153, 153); cursor: default; }

.wvGCSb-PrY1nf .wvGCSb-PLt2Ue-XHP5j:hover { text-decoration: none; }

.wvGCSb-PLt2Ue-QCAl5e { bottom: -10px; color: rgb(17, 85, 204); cursor: pointer; font-size: 12px; padding-right: 5px; padding-top: 5px; position: absolute; right: 5px; text-decoration: none; }

.wvGCSb-PrY1nf .wvGCSb-PLt2Ue-QCAl5e { display: none; }

.wvGCSb-PLt2Ue-I1HBjd { color: rgb(51, 51, 51); padding: 12px 0px 12px 20px; }

.wvGCSb-PLt2Ue-cD65uc { background-color: rgb(254, 247, 224); border-top: 1px solid rgb(218, 220, 224); border-bottom: 1px solid rgb(218, 220, 224); color: rgb(95, 99, 104); font-weight: 500; padding: 12px 20px; position: relative; }

.wvGCSb-PLt2Ue-Q5sUsf, .wvGCSb-PLt2Ue-Q5sUsf:visited { color: rgb(26, 115, 232); font-weight: 400; margin-left: 8px; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-cD65uc { border-top: 0px; box-sizing: border-box; height: 62px; }

.wvGCSb-PLt2Ue-SvJh7b { margin: 6px 29px 10px 20px; position: relative; zoom: 1; }

.wvGCSb-PLt2Ue-SvJh7b-bN97Pc { margin-left: 61px; position: relative; zoom: 1; }

.wvGCSb-PLt2Ue-xqKM5b { font-size: 12px; font-weight: 500; margin-bottom: 3px; top: -3px; }

.wvGCSb-PLt2Ue-r4nke { font-size: 1.2em; margin: 20px 5px 2px; }

.wvGCSb-PLt2Ue-YPqjbf-BeDmAc { top: -4px; }

.wvGCSb-PLt2Ue-YPqjbf-BeDmAc .wvGCSb-YPqjbf-aIWppb { font-weight: 500; }

.wvGCSb-PLt2Ue-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { font-size: 12px; height: 30px; }

.wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(119, 119, 119); line-height: normal; margin-top: 8px; }

.wvGCSb-PLt2Ue-u0pjoe { background-color: rgb(221, 75, 57); border: 1px solid rgb(96, 32, 25); border-radius: 4px; color: rgb(255, 255, 255); margin: 6px; padding: 6px; text-align: center; }

.wvGCSb-PLt2Ue-tJHJj { align-items: center; display: flex; background-color: rgb(245, 245, 245); max-height: 52px; overflow: hidden; padding: 10px 29px 10px 20px; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-tJHJj { background-color: white; border-bottom: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-tJHJj-I5GmGe-ma6Yeb-vFHz9d { border-radius: 8px 8px 0px 0px; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb .HB1eCd-UMrnmb .wvGCSb-PLt2Ue-tJHJj { padding: 12px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-G0jgYd-LgbsSe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-GUUVJe-EnFNjd-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe { margin-right: 4px; width: 40px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe { border-radius: 50%; height: 40px; margin: 0px; padding: 4px; width: 40px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe { line-height: 32px; outline: none; }

.wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { background-color: rgb(232, 234, 237); border: none; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc { top: 5px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { align-items: center; border-radius: 50%; display: flex; height: 32px; justify-content: center; margin: 0px; min-width: 32px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { padding: 4px; }

.wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { display: inline-block; float: left; }

.wvGCSb-F6aDIf .wvGCSb-jNm5if-r4nke-haAclf { align-items: center; display: flex; margin-right: auto; order: -1; }

.wvGCSb-F6aDIf .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS.wvGCSb-jNm5if-tJHJj-r4nke { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 16px; font-weight: 500; line-height: 24px; }

.wvGCSb-PLt2Ue-tJHJj .wvGCSb-yOOK0-EnFNjd { padding: 0px 0px 0px 10px; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-PLt2Ue-tJHJj .wvGCSb-yOOK0-EnFNjd { padding: 0px; width: 160px; }

.wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe { border-color: transparent; background-color: transparent; background-image: none; }

.wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-ZmdkE, .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-auswjd, .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-XpnDCe { border-color: rgb(198, 198, 198); background-color: rgb(248, 248, 248); background-image: -webkit-linear-gradient(top, rgb(248, 248, 248), rgb(241, 241, 241)); }

.wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { visibility: hidden; }

.wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { visibility: visible; }

.wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .wvGCSb-GmVRCe-cHYyed-Bz112c { opacity: 0.3; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-GmVRCe-cHYyed, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GmVRCe-cHYyed { align-items: center; display: flex; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-GmVRCe-cHYyed-Bz112c, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GmVRCe-cHYyed-Bz112c { margin: 0px; }

.wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-OWB6Me .wvGCSb-RmniWd-jNm5if-Bz112c { opacity: 0.15; }

.wvGCSb-PLt2Ue-xxlfEe-haAclf { align-items: center; border-bottom: 1px solid rgb(218, 220, 224); box-sizing: border-box; display: none; justify-content: space-between; max-height: 0px; overflow: hidden; padding: 0px 20px; transition: max-height 0.3s ease-in-out 0s, padding 0.3s ease-in-out 0s; width: 100%; }

.wvGCSb-PLt2Ue-xxlfEe-FNFY6c { display: flex; }

.wvGCSb-PLt2Ue-xxlfEe-PBWx0c { max-height: 100px; padding: 10px 20px; }

.wvGCSb-PLt2Ue-xxlfEe { width: 75%; }

.wvGCSb-PLt2Ue-xxlfEe .wvGCSb-PLt2Ue-G0jgYd-YPqjbf { border: 1px solid rgb(189, 193, 198); border-radius: 8px; box-sizing: border-box; height: auto; padding: 8px 10px; width: 100%; }

.wvGCSb-PLt2Ue-xxlfEe .wvGCSb-PLt2Ue-G0jgYd-YPqjbf:focus { border-color: rgb(77, 144, 254); }

.wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe { margin-right: 8px; }

.wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe-ZmdkE { background-color: transparent; }

.wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { display: none; }

.wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-Bz112c-SxQuSe { width: 18px; height: 18px; margin: 1px 2px 2px 1px; }

.HB1eCd-Bz112c.HB1eCd-HzV7m.wvGCSb-PLt2Ue-GUUVJe-EnFNjd-Bz112c-SxQuSe { width: 24px; height: 24px; margin: 1px 2px 2px 1px; }

.wvGCSb-RXQi4b-HB1eCd-tJHJj .wvGCSb-gkA7Yd-nUpftc { position: relative; overflow: auto; }

.wvGCSb-RXQi4b-HB1eCd-tJHJj .wvGCSb-gkA7Yd-nUpftc-NBtyUd { max-height: 369px; }

.wvGCSb-RXQi4b-HB1eCd-tJHJj:not(.HB1eCd-UMrnmb) .wvGCSb-gkA7Yd-nUpftc > .wvGCSb-dhWRR:first-child { border-top-color: transparent; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-gkA7Yd-nUpftc { bottom: 1px; max-height: none; overflow: hidden auto; position: absolute; top: calc(116px); width: 100%; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-iQd6Fc.wvGCSb-gkA7Yd-nUpftc { margin-top: 40px; }

.HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-gkA7Yd-nUpftc.s4YTVd-NBtyUd-IT5dJd-ORHb { top: calc(170px); }

.wvGCSb-RmniWd-jNm5if-Bz112c { display: inline-block; vertical-align: middle; margin: 4px 5px 5px 2px; opacity: 0.65; }

.HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-Bz112c { opacity: 1; }

.HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-LgbsSe { box-shadow: none; background-color: white; background-image: none; cursor: pointer; border-radius: 2px; border-width: initial; border-style: none; border-image: initial; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; line-height: 16px; padding: 2px 6px 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { background-color: transparent; color: transparent; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { border-radius: 50%; }

.HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { box-shadow: none; background-color: rgb(0, 0, 0); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(241, 243, 244); border-radius: 50%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background-color: rgb(232, 234, 237); border-radius: 50%; }

.HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd { box-shadow: none; background-color: rgb(0, 0, 0); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd { background-color: rgb(232, 234, 237); outline: none; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { align-items: center; font-family: "Google Sans"; font-size: 14px; font-weight: 500; line-height: 28px; text-transform: none; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { align-items: center; color: rgb(60, 64, 67); font-family: "Google Sans"; font-size: 14px; font-weight: 500; line-height: 28px; text-transform: none; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { align-items: center; border: 1px solid rgb(218, 220, 224); border-radius: 24px; color: rgb(95, 99, 104); display: flex; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf { background-color: rgb(232, 240, 254); border: none; color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c-RJLb9c { content: ""; }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c { display: inline-block; margin-bottom: 4px; margin-right: 0px; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae .HB1eCd-Bz112c { display: none; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-cHYyed { margin-left: 4px; }

.HB1eCd-UMrnmb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-cHYyed { overflow: hidden; text-overflow: ellipsis; white-space: nowrap; width: 100px; }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { color: rgb(32, 33, 36); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { color: rgb(24, 90, 188); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { color: rgb(24, 90, 188); background-color: rgb(248, 251, 255); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { background-color: rgb(233, 241, 254); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd { background-color: rgb(225, 236, 254); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { background: rgba(60, 64, 67, 0.04); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { background: rgba(60, 64, 67, 0.12); border: 1px solid rgb(32, 33, 36); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd { background: rgba(60, 64, 67, 0.16); border: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(95, 99, 104); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(26, 115, 232); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(32, 33, 36); }

.HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(24, 90, 188); }

.wvGCSb-yOOK0-EnFNjd-Guievd-WqyaDf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { filter: invert(100%); }

.wvGCSb-yOOK0-EnFNjd-Guievd-WqyaDf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { outline: transparent solid 1px; }

.wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { padding: 2px 0px; }

.HB1eCd-UMrnmb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-OWB6Me { background-color: white; color: rgb(241, 243, 244); cursor: default; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld { cursor: grab; border-color: rgb(232, 234, 237); border-style: solid; border-width: 1px 0px 0px; height: 8px; width: 100%; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld-Bz112c { height: 4px; margin: 2px auto 0px; width: 20px; }

.HB1eCd-UMrnmb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld:hover { background-color: rgb(232, 234, 237); cursor: grab; }

.wvGCSb-PLt2Ue-NkyfNe-imnzkf-m9bMae-MJoBVe-bN97Pc { color: rgb(128, 134, 139); padding-top: 24px; text-align: center; }

.wvGCSb-iQd6Fc .ZYIfFd-IT5dJd-iQd6Fc { display: none !important; }

.ti6hGc-IT5dJd-iQd6Fc { display: none; }

.wvGCSb-iQd6Fc .ti6hGc-IT5dJd-iQd6Fc { display: inline-block !important; }

.wvGCSb-aZ2wEe { height: 100px; overflow: hidden; position: relative; }

.wvGCSb-vyDMJf-aZ2wEe { height: 28px; left: 50%; margin-left: -14px; position: absolute; top: 36px; width: 28px; }

.wvGCSb-vyDMJf-aZ2wEe.auswjd { animation: 1568ms linear 0s infinite normal none running container-rotate; }

.auswjd .aZ2wEe-pbTTYe.aZ2wEe-v3pZbf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running blue-fade-in-out; }

.auswjd .aZ2wEe-pbTTYe.aZ2wEe-oq6NAc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running red-fade-in-out; }

.auswjd .aZ2wEe-pbTTYe.aZ2wEe-gS7Ybc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running yellow-fade-in-out; }

.auswjd .aZ2wEe-pbTTYe.aZ2wEe-nllRtd { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running green-fade-in-out; }

.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running left-spin; }

.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running right-spin; }

.HB1eCd-gkA7Yd-Wz3zdc-haAclf { display: flex; align-items: center; }

.wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-oQLbGe { margin: 0px; }

.wvGCSb-gkA7Yd-Wz3zdc-bN97Pc .wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-oQLbGe .wvGCSb-oQLbGe { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 18px; letter-spacing: 0.25px; line-height: 20px; margin: 0px; max-width: 80%; }

.wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-Wz3zdc { height: 18px; width: 18px; margin-right: 10px; }

.wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-Wz3zdc.wvGCSb-gkA7Yd-Wz3zdc-Wz3zdc-sLO9V-qnnXGd { font-family: "Noto Color Emoji", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 17px; margin-top: -1px; }

.wvGCSb-gkA7Yd-Wz3zdc-bN97Pc { padding-left: 40px; }

.wvGCSb-gkA7Yd-Wz3zdc-tL9eOd { display: flex; }

.wvGCSb-Wz3zdc-nUpftc-YLEF4c { left: 16px; }

.HB1eCd-Hn6s1b { align-items: center; border-radius: 8px; display: flex; flex-direction: row; padding: 12px; }

.HB1eCd-Hn6s1b-Tswv1b { background: rgb(232, 240, 254); }

.HB1eCd-Hn6s1b-Tswv1b > .HB1eCd-Bz112c-RJLb9c { content: ""; }

.HB1eCd-Hn6s1b-lHjamb { background: rgb(254, 239, 195); }

.HB1eCd-Hn6s1b-GMvhG { background: rgb(251, 188, 4); }

.HB1eCd-Hn6s1b-lHjamb > .HB1eCd-Bz112c-RJLb9c, .HB1eCd-Hn6s1b-GMvhG > .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_dark.svg"); }

.HB1eCd-Hn6s1b > .HB1eCd-Bz112c { flex-shrink: 0; height: 24px; width: 24px; }

.HB1eCd-Hn6s1b-Ne3sFf { color: rgb(32, 33, 36); font: 400 14px / 20px Roboto, sans-serif; letter-spacing: 0.2px; margin-left: 12px; }

.wvGCSb-XS83If-suEOdc { display: inline-block; max-width: 35ch; text-align: center; }

.wvGCSb-XS83If-bN97Pc { box-sizing: border-box; text-align: left; width: 330px; }

.wvGCSb-XS83If-bN97Pc.VIpgJd-xl07Ob { border-radius: 8px; white-space: normal; }

.wvGCSb-XS83If-bN97Pc .HB1eCd-Hn6s1b { margin-bottom: 12px; }

.wvGCSb-XS83If-bN97Pc [role="heading"] { color: rgb(32, 33, 36); font: 400 18px / 24px "Google Sans", sans-serif; margin-bottom: 20px; }

.wvGCSb-XS83If-bN97Pc p { color: rgb(95, 99, 104); font: 500 11px / 16px Roboto, sans-serif; letter-spacing: 0.8px; margin-bottom: 16px; text-transform: uppercase; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf { padding: 0px; display: block; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf.tk3N6e-Ru3Ixf-OWB6Me { opacity: 0.38; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf + .tk3N6e-Ru3Ixf { margin-top: 16px; }

.wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-GCYh9b { border: 2px solid rgb(95, 99, 104); height: 15px; width: 15px; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-GCYh9b { left: 3px; top: 50%; transform: translateY(-50%) scale(1.2); }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-ZmdkE:not(.tk3N6e-Ru3Ixf-OWB6Me) .tk3N6e-Ru3Ixf-GCYh9b { cursor: pointer; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-GCYh9b::before { border-color: transparent; border-radius: 50%; border-style: solid; border-width: 6px; content: ""; height: 19px; left: -10.5px; position: absolute; top: -10.5px; transform: scale(0.8333); width: 19px; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc :not(.tk3N6e-Ru3Ixf-OWB6Me):not(.tk3N6e-Ru3Ixf-XpnDCe) .tk3N6e-Ru3Ixf-GCYh9b:hover::before { border-color: rgba(0, 0, 0, 0.06); }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-XpnDCe .tk3N6e-Ru3Ixf-GCYh9b::before { border-color: rgb(232, 240, 254); }

.wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie .tk3N6e-Ru3Ixf-GCYh9b { border-color: rgb(26, 115, 232); }

.wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie.tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-GCYh9b::after { background-color: rgb(26, 115, 232); border-color: rgb(26, 115, 232); border-width: 2px; height: 7px; left: 2px; margin: 0px; top: 2px; width: 7px; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-V67aGc { margin-left: 36px; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-V67aGc label { color: rgb(60, 64, 67); display: block; font: 500 14px / 24px "Google Sans", sans-serif; letter-spacing: 0.1px; }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie .tk3N6e-Ru3Ixf-V67aGc label { color: rgb(26, 115, 232); }

.wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-V67aGc span { color: rgb(95, 99, 104); font: 400 12px / 16px Roboto, sans-serif; letter-spacing: 0.3px; }

.wvGCSb-XS83If-bN97Pc hr { border-right: none; border-bottom: none; border-left: none; border-image: initial; border-top: 1px solid rgb(189, 193, 198); margin: 16px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge .HB1eCd-Bz112c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .EX2EHc-INgbqf-hxXJme-xl07Ob-LgbsSe .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .HB1eCd-Bz112c { height: 18px; width: 18px; margin: 1px 2px 2px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531.svg"); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531.svg"); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-fuEl3d-n9v5ye .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c-haAclf { height: 13220px; position: absolute; width: 83px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-RJLb9c-haAclf { opacity: 0.54; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-RJLb9c-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-OMz1o, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-usbjsf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-EgTfg, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-hDEnYe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-I9GLp, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-nA1mMd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-wlNA0d, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-jSFuyb { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf .HB1eCd-Bz112c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .HB1eCd-Bz112c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge .HB1eCd-Bz112c { margin-top: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c::before, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-dJzjXc-PvRhvb-AznF2e-gk6SMd .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-vOE8Lb-auswjd-AznF2e .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .pD2Zae-Cs2axe-LQ3nce-EfADOe-r4nke .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R.HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-SjW3R-ORHb-Bz112c .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc.HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-F9IAbd-HSrbLb-JMoATd.HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-NkY1gc-fFW7wc-LgbsSe-nVMfcd .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .F9IAbd-UzWXSb-gElRsf-MZArnb-VCkuzd-pIkB8-qAJZhe-LgbsSe .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .Td0Hgc-YjoMNe-VCkuzd-v3pZbf-Bz112c .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec .HB1eCd-Bz112c-RJLb9c, .HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.lUepf-nEeMgc .HB1eCd-Bz112c { margin: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-QbdDtf-oKdM2c-Bz112c .RbRzK-Bz112c { margin: -1px 0px 0px -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-sLO9V-rdwzAe { font-family: "Google Symbols"; height: 0px; position: absolute; overflow: hidden; width: 0px; z-index: -1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-w7bdYb-iyXyEd { left: 0px; top: -9674px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Q4BLdf { left: 0px; top: -9014px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-jNm5if { left: -40px; top: -7146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-HB1eCd { left: 0px; top: -11530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-RFAvhb { left: 0px; top: -11838px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-Va8Ffe-a1e4Ad { left: 0px; top: -2826px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-iyXyEd { left: 0px; top: -11818px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-xJzy8c { left: 0px; top: -9164px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-htvI8d-wcotoc-ndfHFb { left: -40px; top: -1438px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-cGMI2b { left: -40px; top: -3060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-oXtfBe { left: -60px; top: -3060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-oXtfBe { left: -20px; top: -8792px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-LK5yu { left: -26px; top: -7890px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-DKlKme-qwU8Me { left: -20px; top: -12210px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-yIbDgf { left: 0px; top: -2356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-LK5yu { left: 0px; top: -6876px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-AipIyc { left: 0px; top: -4020px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-qwU8Me { left: 0px; top: -12506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-ma6Yeb { left: -42px; top: -8690px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-cGMI2b { left: -48px; top: -13172px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-oXtfBe { left: -26px; top: -7646px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fW01td-BvBYQ-ma6Yeb { left: -40px; top: -3102px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XXCpLd-Bpn8Yb { left: -62px; top: -11344px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XXCpLd-Bpn8Yb-mlk5z { left: -40px; top: -2978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-OiiCO { left: -22px; top: -11304px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KmuGVc-MHYjYb { left: -52px; top: -10648px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MqcBrc-s4vhY { left: -42px; top: -8730px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-IyROMc-wlNA0d { left: -40px; top: -10466px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o { left: -26px; top: -10012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o-v3pZbf { left: -20px; top: -76px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BoKuKe-OMz1o-MFS4be { left: 0px; top: -2958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XHgP6b-SDqDXe-iAqvw { left: -62px; top: -3472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-XHgP6b-f4z2Dd-E4ZlWe { left: -60px; top: -5388px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-elBQIf { left: -62px; top: -4964px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-c8csvc { left: -20px; top: -3594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-K0TrJc { left: -62px; top: -12668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-HrRdod-yLHjwb { left: -62px; top: -9634px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-km6h5c { left: 0px; top: -4882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QLEXN { left: -42px; top: -1062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QLEXN-DKlKme { left: -42px; top: -5708px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-WPi0i-MR5Q1e { left: 0px; top: -4964px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MPu53c { left: -26px; top: -10222px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-OVkoRd-GEUYHe { left: -15px; top: -484px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JbbQac-Wxxdob { left: 0px; top: -7532px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TvD9Pc { left: 0px; top: -1084px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nyE0bc { left: -42px; top: -1230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-J5uZjd-edvN0e { left: -42px; top: -8770px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-DyVDA { left: 0px; top: -5166px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-DyVDA-mPlZac { left: 0px; top: -11346px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-N7Eqid-GMvhG { left: 0px; top: -608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jNm5if-MCEKJb { left: -22px; top: -11654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bKkSne-obrOwb { left: -26px; top: -10182px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bN97Pc-jCCvxc { left: -42px; top: -3472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-bMcfAe-pKrx3d-lbYRR { left: -26px; top: -1014px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QdThLb { left: -60px; top: -12820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-UkZFS { left: -62px; top: -11304px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xceQUb { left: -20px; top: -8536px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-VkLyEc-zM6fo { left: -20px; top: -5388px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-FuIHKe-R1gDOc-MR5Q1e { left: -40px; top: -6168px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Oo0NPd { left: 0px; top: -3100px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uG5Yqe-JPn0pf-DKlKme { left: -20px; top: -9932px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uG5Yqe-JPn0pf-BvBYQ { left: 0px; top: -5086px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nupQLb { left: -20px; top: -11530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nupQLb-Q4BLdf { left: 0px; top: -2482px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-cXXICe-x5cW0b { left: -42px; top: -8710px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn { left: 0px; top: -7512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn-MFS4be { left: -60px; top: -2114px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-QymXn-oq6NAc { left: 0px; top: -12210px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ndfHFb-aTv5jf { left: 0px; top: -4546px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-j4gsHd-hFsbo-bEDTcc-LkdAo { left: 0px; top: -4040px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DyVDA-D5MPn { left: -20px; top: -12360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DyVDA-D5MPn-ImBhed { left: -26px; top: -8624px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xvr5H-i5vt6e { left: 0px; top: -3182px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wz3zdc { left: -62px; top: -1230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DJPBic-AFZkUd { left: -20px; top: -3684px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fHSeKd-LkdAo { left: -26px; top: -6230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-vgRlPd-XigvTc-rDoBzb { left: 0px; top: -1062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KoToPc { left: -40px; top: -8792px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KoToPc-DKlKme { left: -40px; top: -9932px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hdBvUb { left: 0px; top: -6654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PlOyMe-vOE8Lb-jCCvxc { left: 0px; top: -3532px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TZk80d-ZGNLv-I9GLp { left: -20px; top: -12918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TZk80d-jCCvxc { left: 0px; top: -6586px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-HTFGIc { left: 0px; top: -12002px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-bRSSXe { left: 0px; top: -2868px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-bRSSXe-Hyc8Sd { left: -20px; top: -2754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yOOK0-jyrRxf-nUpftc { left: -20px; top: -1698px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-lCdvJf-bEDTcc-DARUcf { left: 0px; top: -10648px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-lCdvJf-BIr6Bc { left: -20px; top: -3882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-drxrmf-wcotoc-jirZld { left: -62px; top: -11798px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-AHmuwe-oXtfBe { left: -20px; top: -3102px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yEEHq { left: -20px; top: -6028px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-yEEHq-x5cW0b { left: -62px; top: -8150px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-JNdkSc { left: 0px; top: -13074px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-JPn0pf { left: -34px; top: -5926px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Wxxdob-xSQTrd { left: 0px; top: -7444px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sLO9V-fmcmS-SxQuSe { left: -40px; top: -11738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xRdasc-oKdM2c-dJDgTb { left: 0px; top: -4422px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n9oEIb { left: -44px; top: -8812px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n9oEIb-SNIJTd { left: -42px; top: -1738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TBCoIc { left: 0px; top: -3122px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ObfsIf-KzxUkd { left: -42px; top: -12688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ObfsIf-vhhrIe { left: -40px; top: -5514px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-tJHJj-yePe5c { left: -26px; top: -6520px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-h9d3hd { left: -60px; top: -1498px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ZYIfFd-fbudBf { left: -60px; top: -2774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ntN8G { left: 0px; top: -5648px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TIHSC-E8fGCc { left: -52px; top: -8878px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DKlKme-RWgCYc { left: 0px; top: -3320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DKlKme-YMi5E { left: -20px; top: -5608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xguqbd { left: 0px; top: -10668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-YRhSCb { left: 0px; top: -1564px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-YRhSCb-SIsrTd { left: -62px; top: -5660px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-nGOfy { left: -42px; top: -12042px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BKD3ld-nGOfy-SIsrTd { left: -22px; top: -10716px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Tswv1b { left: -20px; top: -10472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-kWbB0e-D5MPn { left: -20px; top: -3554px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-YPqjbf { left: 0px; top: -12400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rYk4U { left: -42px; top: -4712px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-c53jI-TBCoIc { left: -20px; top: -8858px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-O807Gb { left: -60px; top: -8858px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-LIMNJb { left: 0px; top: -320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-LIMNJb-AznF2e { left: 0px; top: -232px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-V67aGc { left: -62px; top: -7512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-mSEUvf { left: -52px; top: -9118px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-QLEXN-VMPhoe { left: -62px; top: -6762px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-wwuYjd { left: -20px; top: -7126px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RWgCYc-yY4Wcc { left: -20px; top: -2114px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd { left: -60px; top: -3882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd-Q4BLdf { left: -62px; top: -3280px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hSRGPd-Xhs9z { left: -62px; top: -5708px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Jn51gd { left: -40px; top: -8476px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Jn51gd-SIsrTd { left: 0px; top: -5388px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rymPhb-Rv62Se { left: -42px; top: -4628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pGuBYc-TvD9Pc { left: -62px; top: -6742px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pGuBYc-FNFY6c { left: -20px; top: -10758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-l4eHX-t02dhe { left: 0px; top: -8750px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JtB1fc { left: -52px; top: -7404px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xSh02c { left: -20px; top: -10506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-H1aTHf { left: -42px; top: -10310px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DUGJie-Q4BLdf { left: 0px; top: -3574px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-z5C9Gb-zcdHbf-BvBYQ { left: 0px; top: -4146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-x5cW0b-nKQ6qf-hgHJW { left: -40px; top: -4292px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-x5cW0b-nKQ6qf-yHKmmc { left: -42px; top: -7512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-h1U9Be { left: 0px; top: -7424px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RFnRab-MCEKJb { left: -60px; top: -9320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-b3rLgd-HzFBSb { left: -20px; top: -2336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Vgu1H-mKZypf { left: -22px; top: -1738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n5AaSd-u3Agqb { left: 0px; top: -1800px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PrY1nf-nQ1Faf { left: -60px; top: -9400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PrY1nf-nQ1Faf-MFS4be { left: -40px; top: -10958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-pBztBd-dJfz0c-JZnCve { left: -40px; top: -12102px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-G84jIc { left: -62px; top: -3842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-FNFY6c-RmniWd-uJ3wk { left: -62px; top: -3662px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-LhcNjd { left: -22px; top: -12022px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-ij8cu { left: 0px; top: -5514px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DARUcf-Lr2Z8d { left: 0px; top: -2436px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RF62N-nEeMgc-Ia7Qfc { left: 0px; top: -10472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KNM5Ef { left: -20px; top: -6210px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-KNM5Ef-Q4BLdf { left: -40px; top: -212px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-g7W7Ed-qwU8Me-wcotoc-LK5yu { left: 0px; top: -170px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Ft5J4b { left: -62px; top: -4984px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Ft5J4b-di8rgd-Wxxdob { left: 0px; top: -9932px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-GEUYHe-JNdkSc { left: -26px; top: -7032px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Faem2b-cVFi4 { left: -48px; top: -8572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-iyXyEd { left: -48px; top: -1014px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-iyXyEd-g6cJHd { left: 0px; top: -11264px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nQ1Faf { left: -22px; top: -3202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nQ1Faf-Xhs9z { left: -26px; top: -9538px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xJzy8c-HiaYvf { left: -44px; top: -4400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xJzy8c-HiaYvf-O1htCb { left: 0px; top: -12420px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Jz7rA { left: 0px; top: -980px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-zSI2l-QLEXN { left: 0px; top: -6168px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-n8nH7-jyrRxf { left: 0px; top: -9206px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jRmmHf-ibnC6b { left: -20px; top: -6676px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NziyQe-LkdAo { left: -52px; top: -6518px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TdyTDe { left: -20px; top: -5688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-TdyTDe-r9oPif { left: 0px; top: -9138px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-g3I98d { left: 0px; top: -2242px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-aIWppb-htvI8d { left: -46px; top: -5044px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EgTfg { left: -40px; top: -3554px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EgTfg-gS7Ybc { left: -40px; top: -2876px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PEFSMe { left: 0px; top: -9320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-xXq91c-oQYOj { left: 0px; top: -4292px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Gpz5id { left: -40px; top: -8858px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-uXLMpd { left: -60px; top: -8536px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qrlFte { left: -22px; top: -11674px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Iqlsrf { left: -58px; top: -6068px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-S9gUrf-HiaYvf { left: -60px; top: -10486px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-m3mY0d-Q4BLdf { left: 0px; top: -12380px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qwU8Me-rrhWne { left: 0px; top: -8792px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ReqAjb-qwU8Me-MnhZ9d { left: 0px; top: -8834px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-ktSouf { left: -40px; top: -12820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NgtDm-YS35zb { left: -54px; top: -5004px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-O1htCb-NkyfNe { left: -20px; top: -11490px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EnFNjd-ryxqyc { left: -40px; top: -2814px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JPn0pf { left: 0px; top: -10248px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RFAvhb-AznF2e { left: -26px; top: -2502px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-if5aCc-sTBVle { left: -42px; top: -11674px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-luNtDf-s2ctBd { left: 0px; top: -13116px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-V5oUn { left: -20px; top: -2868px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb { left: -60px; top: -10506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb-e7aFhf { left: -20px; top: -1438px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Bpn8Yb-uTrtOd { left: -40px; top: -2336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-rvOPdc-RFnRab { left: 0px; top: -300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-JK9eJ { left: 0px; top: -8496px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DIdRlc { left: -40px; top: -11510px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-DIdRlc-nyE0bc { left: 0px; top: -8690px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hDEnYe-JaPV2b { left: -22px; top: -2548px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-hDEnYe-nllRtd { left: 0px; top: -5668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-Q4BLdf-gvZm2b { left: -20px; top: -608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-ObfsIf-nUpftc { left: 0px; top: -8476px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BaYisc-uaxL4e { left: -62px; top: -1130px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i2RYZ { left: 0px; top: -192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sTBVle-BvBYQ { left: -52px; top: -7424px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Yygnk { left: -42px; top: -11404px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Yygnk-Z5I80b { left: -26px; top: -7672px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-QLEXN { left: -60px; top: -6296px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-g6cJHd { left: -40px; top: -11550px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-jyrRxf-AznF2e { left: -42px; top: -11654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-sAb8f { left: -60px; top: -3902px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-rrhWne-hgHJW { left: -20px; top: -5988px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-rrhWne-yHKmmc { left: -20px; top: -9952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-hgHJW { left: 0px; top: -5146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-tSZMSb { left: 0px; top: -3902px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-yHKmmc { left: -20px; top: -6190px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-fmcmS-ReqAjb-BvBYQ-EbqdBd { left: -60px; top: -3080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-EWK8Bb { left: -20px; top: -2958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-RCfa3e { left: -62px; top: -252px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-L4Nn5e { left: -20px; top: -11940px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-e3BBL-yHKmmc-hFsbo { left: -20px; top: -11510px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-Zj4Smb-Z5I80b-GMvhG { left: 0px; top: -1020px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-NowJzb { left: 0px; top: -6316px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-sfGayb { left: -42px; top: -11818px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-MHYjYb-J6RZ7b { left: -40px; top: -8750px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-zf3vf { left: 0px; top: -3594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-dIxMhd-DyVDA-TIHSC { left: 0px; top: -6008px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-dIxMhd-iWMRLe-EnFNjd { left: 0px; top: -11570px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-BvBYQ-nyE0bc { left: -46px; top: -12460px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nUpftc-kPTQic { left: -60px; top: -2436px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nUpftc-ti6hGc { left: -22px; top: -2896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-qPaVXd-yHKmmc { left: 0px; top: -212px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-PJVNOc-hYO5Oc { left: -42px; top: -8670px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-ltEGzf { left: 0px; top: -8858px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-RPzgNd { left: 0px; top: -4822px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-i8xkGf-fmcmS-i8xkGf { left: -40px; top: -12230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-nJjxad-bEDTcc { left: -58px; top: -5278px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-h30Snd-ovCUCd { left: -42px; top: -12002px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-h30Snd-ovCUCd-r9oPif { left: -46px; top: -9206px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb-ovCUCd { left: 0px; top: -340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ktSouf { left: -60px; top: -2978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PEFSMe { left: -60px; top: -12506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PEFSMe-E3DyYd { left: -20px; top: -1252px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-SIsrTd { left: -40px; top: -6028px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-E3DyYd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-SIsrTd-E3DyYd { left: -20px; top: -8670px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-SIsrTd { left: 0px; top: -6546px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uXLMpd-E3DyYd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-SIsrTd-E3DyYd { left: -58px; top: -2592px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc { left: 0px; top: -12820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc-r9oPif { left: -26px; top: -4080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-UkZFS { left: 0px; top: -11510px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b { left: -60px; top: -12860px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-OMz1o { left: 0px; top: -11408px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EgTfg, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-usbjsf { left: -20px; top: -2436px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EgTfg-TLxrU { left: 0px; top: -11124px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hDEnYe { left: -60px; top: -9300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-I9GLp { left: 0px; top: -10268px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-I9GLp-JaPV2b { left: -60px; top: -6276px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd { left: -52px; top: -4754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jSFuyb { left: -40px; top: -9300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd-JaPV2b { left: 0px; top: -1458px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nA1mMd-JaPV2b-r9oPif { left: -40px; top: -5682px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TFrYib { left: -40px; top: -11880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-oO2eQ { left: 0px; top: -2628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PJVNOc { left: 0px; top: -10758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-wlNA0d { left: 0px; top: -3040px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-wlNA0d { left: -20px; top: -7444px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jbwjpc-RvIlWb { left: -52px; top: -9834px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lcE6r-JLm1tf-YZ04zc-RvIlWb { left: -52px; top: -4566px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-N7Eqid-RvIlWb { left: 0px; top: -8218px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-Xhs9z-RvIlWb { left: 0px; top: -5900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vVQOP { left: -40px; top: -7356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-AV3gEe-Q4BLdf-XpSwdc { left: 0px; top: -10426px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf { left: -48px; top: -1034px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eFD6re { left: 0px; top: -6722px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-c8csvc { left: -20px; top: -668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-c8csvc-E3DyYd { left: 0px; top: -6632px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-O807Gb { left: -62px; top: -9786px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-O807Gb-E3DyYd { left: -22px; top: -11716px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-hxXJme { left: -40px; top: -1458px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-hxXJme-E3DyYd { left: 0px; top: -2528px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-LK5yu { left: -62px; top: -6830px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-LK5yu-E3DyYd { left: 0px; top: -9538px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-oXtfBe { left: -40px; top: -2958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-oXtfBe-E3DyYd { left: -20px; top: -2072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-qwU8Me { left: -20px; top: -2978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-qwU8Me-E3DyYd { left: -20px; top: -3512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-yIbDgf { left: -62px; top: -12918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-yIbDgf-E3DyYd { left: 0px; top: -11980px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-LK5yu { left: -48px; top: -1938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-oXtfBe { left: 0px; top: -7356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-qwU8Me { left: -52px; top: -11084px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-ma6Yeb { left: 0px; top: -7124px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-AipIyc { left: -20px; top: -8650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fW01td-JPn0pf-cGMI2b { left: -60px; top: -9932px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uG5Yqe-JPn0pf-agdLee { left: 0px; top: -1872px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uG5Yqe-JPn0pf-o7abwc { left: -40px; top: -6190px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-ma6Yeb { left: 0px; top: -12572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-ma6Yeb-E3DyYd { left: 0px; top: -9054px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-AipIyc { left: 0px; top: -10938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-AipIyc-E3DyYd { left: 0px; top: -6402px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-cGMI2b { left: 0px; top: -1438px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tHaKme-cGMI2b-E3DyYd { left: -26px; top: -7592px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H { left: -26px; top: -6588px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-E3DyYd { left: 0px; top: -4712px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-r9oPif { left: -48px; top: -1370px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Rv62Se-EXHrde-Ca4zAd { left: 0px; top: -6424px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv { left: 0px; top: -11758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-E3DyYd { left: -60px; top: -5470px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-r9oPif { left: -20px; top: -12400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Jn51gd-EXHrde-Ca4zAd { left: -22px; top: -2722px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld { left: -26px; top: -9482px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-E3DyYd { left: -20px; top: -6456px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc { left: 0px; top: -6742px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-E3DyYd { left: -46px; top: -6230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd { left: 0px; top: -1000px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-E3DyYd { left: -46px; top: -5064px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nyE0bc { left: -20px; top: -11798px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NowJzb { left: -62px; top: -1110px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NowJzb-E3DyYd { left: -36px; top: -170px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-yTCTk { left: -20px; top: -3534px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-I7wDP { left: -48px; top: -7772px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-I7wDP-r9oPif-T60B1 { left: 0px; top: -12460px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf { left: 0px; top: -10918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf-E3DyYd { left: -52px; top: -5900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JPn0pf-r9oPif-gS7Ybc { left: -26px; top: -582px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .EX2EHc-Bz112c-LSk3jc-BHsdwc { left: 0px; top: -10114px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QBLLGd { left: -55px; top: -5112px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-weuhHc-E3DyYd { left: -48px; top: -9254px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-FXrc0c { left: 0px; top: -6190px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-wZVHld-V67aGc { left: -52px; top: -6696px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tJiF1e { left: 0px; top: -3362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MYFTse { left: -22px; top: -6916px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-di8rgd-hxXJme { left: 0px; top: -6230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-edvN0e-hxXJme { left: -60px; top: -2918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-edvN0e-hxXJme-E3DyYd { left: -26px; top: -3018px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-hxXJme { left: -40px; top: -3902px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-rTEl { left: -20px; top: -11694px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-SX9D7d-E3DyYd { left: 0px; top: -3842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf { left: -40px; top: -6722px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-r9oPif { left: 0px; top: -7572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-nUpftc-ZdbLkb { left: -60px; top: -9054px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-eKpHRd-BPrWId-r9oPif { left: -46px; top: -11224px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if { left: -42px; top: -9676px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-jNm5if-E3DyYd { left: -52px; top: -8594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e { left: -20px; top: -3122px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-E3DyYd { left: -48px; top: -13094px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-AHUcCb { left: -60px; top: -4060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-E3Uge { left: -20px; top: -1498px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-Qs3R8d-E3DyYd { left: -60px; top: -7356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-J2Tr8e-uPjwvb-ZdbLkb { left: -42px; top: -12572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-jNm5if { left: -20px; top: -2242px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-jNm5if-r9oPif { left: 0px; top: -2774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-yHKmmc-r9oPif { left: -48px; top: -12184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-yHKmmc-yaNpec { left: 0px; top: -9744px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e3BBL-hgHJW-yaNpec { left: 0px; top: -7336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QLEXN { left: -20px; top: -3162px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-QLEXN-E3DyYd { left: -42px; top: -6916px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QLEXN-r9oPif { left: -48px; top: -7572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-SIsrTd { left: -22px; top: -8770px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-Vgu1H-SIsrTd-E3DyYd { left: -52px; top: -3382px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-SIsrTd { left: -62px; top: -11384px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-ZGNLv-SIsrTd-E3DyYd { left: -60px; top: -11940px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-SIsrTd { left: -60px; top: -8750px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-BKD3ld-SIsrTd-E3DyYd { left: -20px; top: -9744px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-SIsrTd { left: 0px; top: -4842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-CYXvYc-SIsrTd-E3DyYd { left: -26px; top: -9254px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-SIsrTd { left: 0px; top: -5106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-wwuYjd-SIsrTd-E3DyYd { left: -42px; top: -1252px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-i3jM8c { left: -22px; top: -9676px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-i3jM8c-E3DyYd { left: -60px; top: -9952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-SIsrTd { left: -40px; top: -11530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-SIsrTd-E3DyYd { left: -60px; top: -6168px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vOE8Lb-SIsrTd { left: 0px; top: -11244px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vOE8Lb-SIsrTd-E3DyYd { left: -44px; top: -10978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf { left: 0px; top: -862px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LQY1ye { left: -62px; top: -11858px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zjQX3e { left: -62px; top: -4692px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i2RYZ { left: -60px; top: -3554px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i2RYZ-E3DyYd { left: 0px; top: -11284px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JbbQac-TCl01b { left: -20px; top: -5514px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd { left: -40px; top: -1498px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-E3DyYd { left: 0px; top: -7166px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-dJfz0c-JZnCve { left: -42px; top: -3300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-dJfz0c-JZnCve-r9oPif { left: -56px; top: -5952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-HLvlvd { left: -42px; top: -11304px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-purZT { left: 0px; top: -668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-SdkFre { left: 0px; top: -1758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RF62N-Wxxdob { left: -20px; top: -11738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RF62N-Wxxdob-E3DyYd { left: -20px; top: -11570px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf { left: -52px; top: -7444px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL { left: -40px; top: -12062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL-SIsrTd { left: 0px; top: -2754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DARUcf-LhcNjd { left: -22px; top: -12042px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DARUcf-LhcNjd-r9oPif { left: -22px; top: -13120px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc { left: 0px; top: -1658px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd { left: -62px; top: -9766px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yHKmmc { left: 0px; top: -1892px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hgHJW { left: 0px; top: -5608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-DARUcf { left: -48px; top: -9718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xvr5H { left: -20px; top: -3492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vgRlPd { left: -48px; top: -1918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vgRlPd-r9oPif { left: 0px; top: -2046px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DKlKme-RWgCYc { left: 0px; top: -3684px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-DKlKme-RWgCYc-r9oPif { left: 0px; top: -3778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-oXtfBe-VBrcT { left: -22px; top: -4712px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-oXtfBe-cGMI2b-VBrcT { left: -60px; top: -2754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-LK5yu-VBrcT { left: -20px; top: -628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-R8Knhb-qwU8Me-VBrcT { left: -42px; top: -2072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mQXP-r9oPif { left: -40px; top: -5634px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-CtVXDf-r08add-BKD3ld-cXXICe-VBrcT { left: -26px; top: -9472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-NkyfNe { left: -62px; top: -10248px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-NkyfNe-E3DyYd { left: -46px; top: -1084px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-qwU8Me { left: 0px; top: -7146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-qwU8Me-E3DyYd { left: -22px; top: -4942px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-LK5yu { left: 0px; top: -6856px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-LK5yu-E3DyYd { left: -48px; top: -1820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-ma6Yeb { left: -26px; top: -9906px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-ma6Yeb-E3DyYd { left: -22px; top: -11980px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-cGMI2b { left: 0px; top: -12918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-cGMI2b-E3DyYd { left: -52px; top: -4774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-sfSLhd { left: 0px; top: -4166px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-sfSLhd-E3DyYd { left: -48px; top: -9608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-EcYfVc { left: -20px; top: -9184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-EcYfVc-E3DyYd { left: -48px; top: -8432px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-tSZMSb { left: 0px; top: -11694px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-tSZMSb-E3DyYd { left: -20px; top: -10526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-DKlKme { left: -62px; top: -8770px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-DKlKme-E3DyYd { left: 0px; top: -6498px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-BvBYQ { left: -62px; top: -11878px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-BvBYQ-E3DyYd { left: 0px; top: -6916px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xSh02c { left: -20px; top: -2826px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf { left: -40px; top: -12210px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd { left: -26px; top: -12460px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pXHOFf { left: 0px; top: -5024px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pXHOFf-MFS4be { left: -20px; top: -4060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-s2ctBd { left: -26px; top: -556px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-s2ctBd-E3DyYd { left: -52px; top: -2154px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-NUaK6d { left: -20px; top: -1892px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-PoC6nf { left: -46px; top: -7890px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-PoC6nf-i5vt6e { left: -44px; top: -7910px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e { left: -20px; top: -12526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e-ZmdkE { left: -22px; top: -1718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-i5vt6e-QDgCrf { left: 0px; top: -5628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-Hyc8Sd { left: 0px; top: -9184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb { left: -52px; top: -9492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-LkdAo-r9oPif { left: 0px; top: -7844px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-hJDwNd { left: 0px; top: -38px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-hJDwNd-sM5MNb { width: 36px; height: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-a4fUwd { left: -60px; top: -8792px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-a4fUwd-SIsrTd { left: -60px; top: -11510px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-z5C9Gb { left: -26px; top: -3804px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-z5C9Gb-SIsrTd { left: 0px; top: -11880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-UlV2sd-OMz1o { left: -42px; top: -1758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-uPjwvb { left: -26px; top: -9808px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-h0Nkge-uPjwvb-r9oPif { left: 0px; top: -3804px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qrlFte-uPjwvb-r9oPif { left: -48px; top: -9880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd { left: -48px; top: -12142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-E3Uge { left: 0px; top: -11798px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-NkyfNe { left: -48px; top: -1418px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PJVNOc-hYO5Oc { left: 0px; top: -12082px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-PvhD9 { left: 0px; top: -2938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ij8cu-r9oPif { left: -52px; top: -11592px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd { left: -20px; top: -11960px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe { left: 0px; top: -5688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe-HLvlvd { left: -60px; top: -8476px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-O0r3Gd { left: -40px; top: -1564px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-O0r3Gd-u0pjoe-r9oPif-Qhstab { left: -20px; top: -4822px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zM6fo { left: -22px; top: -1758px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8 { left: -40px; top: -6362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8-E3Uge { left: 0px; top: -7870px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pmuK7 { left: 0px; top: -7104px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-fZiSAe { left: -42px; top: -9786px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pX1iqf-kPTQic { left: -40px; top: -6830px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-SNIJTd-kPTQic { left: 0px; top: -5126px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-DyVDA { left: 0px; top: -11940px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-DyVDA-ImBhed { left: -26px; top: -4800px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-nUpftc { left: -60px; top: -2336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd { left: -26px; top: -9144px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-VCkuzd-TLxrU { left: 0px; top: -6456px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-VCkuzd-HLvlvd { left: -42px; top: -12918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-iyXyEd-TLxrU { left: 0px; top: -10958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l03kKd-iyXyEd-JH1xTd-TLxrU { left: -20px; top: -3142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd-htvI8d-HLvlvd { left: -26px; top: -6628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc { left: -22px; top: -12688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lbYRR { left: 0px; top: -842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d { left: -42px; top: -10072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G84jIc { left: 0px; top: -7012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-V67aGc-S8vSze { left: 0px; top: -4692px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pKrx3d-SxQuSe { left: -60px; top: -10526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xXq91c { left: 0px; top: -7378px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-T3yXSc { left: 0px; top: -12840px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-BvBYQ-kolMJb { left: -42px; top: -12708px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LK5yu-kqOKYb { left: -62px; top: -8670px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qwU8Me-kqOKYb { left: 0px; top: -12062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LK5yu-kqOKYb-kolMJb { left: -20px; top: -9320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qwU8Me-kqOKYb-kolMJb { left: 0px; top: -12800px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf { left: -20px; top: -4292px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-x5cW0b { left: -20px; top: -3902px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DltcQc-CCJ0ld { left: -22px; top: -4732px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NMrWyd-s3Bhse { left: -52px; top: -8218px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hj4D6d-vJ7A6b { left: -60px; top: -1658px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-bEDTcc-E3DyYd { left: -20px; top: -1062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-m9bMae { left: -26px; top: -8078px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-yY4Wcc { left: -62px; top: -4628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nupQLb { left: 0px; top: -6676px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MrxDPd-jyrRxf { left: 0px; top: -1110px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hDEnYe-jkpPIb { left: 0px; top: -11920px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-Q9HdGd { left: -20px; top: -4106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QbShld { left: 0px; top: -6382px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zcdHbf { left: 0px; top: -12122px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sJY2Bf-bVEB4e { left: -40px; top: -3492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf { left: 0px; top: -6566px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-OiiCO { left: -40px; top: -3882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-r9oPif { left: 0px; top: -530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-u0pjoe-u2z5K { left: -42px; top: -2180px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sKFHqe { left: -20px; top: -13074px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sKFHqe-SIsrTd { left: -20px; top: -6168px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NBDE7b { left: -46px; top: -3822px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod { left: -60px; top: -2794px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-CBeBSd-EFlEBf { left: 0px; top: -9634px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-VgwJlc-xTMeO { left: -20px; top: -4964px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-VgwJlc-FNFY6c { left: -60px; top: -608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc { left: -20px; top: -4984px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc-r9oPif { left: -48px; top: -2998px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ud7fr { left: -20px; top: -11880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-R1s0ee-uDEFge-yaNpec { left: 0px; top: -816px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ud7fr-r9oPif { left: -20px; top: -10622px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-v3pZbf { left: -62px; top: -3300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-aVTXAb { left: -40px; top: -2754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sI3MNd { left: -52px; top: -12754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed { left: -52px; top: -10710px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-E3DyYd { left: -52px; top: -10688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-K0TrJc-JaPV2b { left: -26px; top: -2998px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-aVTXAb-v3pZbf { left: -60px; top: -9360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc { left: -62px; top: -10132px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c { left: -62px; top: -10288px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c-rTEl { left: -40px; top: -4106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-rTEl { left: -26px; top: -6608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-rTEl { left: 0px; top: -4902px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl { left: -40px; top: -4146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl-E3DyYd { left: -52px; top: -9564px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-rTEl-r9oPif { left: -48px; top: -7078px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GCYh9b-rTEl { left: -46px; top: -816px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-skjTt-rTEl { left: -40px; top: -9320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-rTEl { left: 0px; top: -3080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ihIZgd-rTEl { left: -26px; top: -7572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-r9oPif { left: -56px; top: -6382px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-fmcmS-eEGnhe { left: -22px; top: -6402px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-IT5dJd { left: 0px; top: -7798px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-IT5dJd-HLvlvd { left: -62px; top: -4822px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EXxX1b-Q9HdGd-Xhs9z { left: -26px; top: -4334px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-nGOfy { left: -52px; top: -12552px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-nGOfy-E3DyYd { left: 0px; top: -1348px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-YRhSCb { left: 0px; top: -10526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cjo6sd-YRhSCb-E3DyYd { left: 0px; top: -4922px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-HLvlvd { left: -52px; top: -11042px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-di8rgd-YwNhXd { left: -22px; top: -4692px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QdThLb { left: -42px; top: -10052px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QdThLb-E3DyYd { left: 0px; top: -2846px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nllRtd-g6cJHd { left: -42px; top: -4250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sLO9V-SxQuSe { left: -52px; top: -10668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf-HiaYvf { left: -20px; top: -10918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-S9gUrf-HiaYvf-E3DyYd { left: 0px; top: -9608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YIAiIb-rDoBzb { left: -60px; top: -4106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Fq92xe-mU4ghb { left: -22px; top: -9634px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yUKnc { left: 0px; top: -2978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-RPzgNd { left: -56px; top: -6408px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-i8xkGf { left: 0px; top: -2134px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i8xkGf-ltEGzf { left: 0px; top: -2092px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-b58pU { left: -62px; top: -11818px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nllRtd-a4fUwd { left: -20px; top: -11346px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-HLvlvd { left: -26px; top: -3228px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-HLvlvd-SIsrTd { left: 0px; top: -9808px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-h9d3hd { left: -20px; top: -5470px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sn54Q-nllRtd { left: -52px; top: -8918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eNZ9Nb { left: -26px; top: -7614px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-r9oPif { left: -46px; top: -9906px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-JaPV2b { left: -60px; top: -2876px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-JaPV2b-nNtqDd { left: -40px; top: -2794px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-nllRtd { left: -20px; top: -1544px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hdBvUb-HLvlvd { left: -22px; top: -11324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-OpAKde-QLEXN { left: -20px; top: -12062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-OpAKde-QLEXN-HLvlvd { left: -22px; top: -4922px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nJjxad-bEDTcc { left: -22px; top: -7166px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc { left: -60px; top: -3100px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc-i5vt6e-J9pn5c-r9oPif { left: -52px; top: -4592px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW { left: -44px; top: -11980px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW-i5vt6e-J9pn5c-r9oPif { left: 0px; top: -9560px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jsmBPd-GMvhG { left: -26px; top: -2482px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KsV2dd { left: -62px; top: -10052px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb { left: 0px; top: -6048px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-B1neQd-TCl01b { left: -40px; top: -9184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-UmQjBf { left: -20px; top: -6742px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-QLEXN { left: -58px; top: -5298px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-to915 { left: -26px; top: -9558px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-qwU8Me-IFdKyd-HLvlvd-r9oPif { left: -52px; top: -10896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-a4fUwd-to915-SIsrTd { left: -46px; top: -2396px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc { left: -52px; top: -10156px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-E3DyYd { left: -20px; top: -10312px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-r9oPif { left: -52px; top: -10176px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-N2TEqe { left: -42px; top: -9766px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ZMv3u-QLEXN { left: 0px; top: -12898px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ZMv3u-QLEXN-i5vt6e-r9oPif { left: -26px; top: -6336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-dJDgTb-QLEXN { left: -62px; top: -10072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-dJDgTb-QLEXN-i5vt6e-r9oPif { left: -26px; top: -6562px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QLEXN { left: -62px; top: -11324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-QLEXN-r9oPif { left: -44px; top: -4922px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN { left: -22px; top: -1230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN-i5vt6e { height: 18px; left: 0px; top: -10288px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zSI2l-QLEXN-i5vt6e-r9oPif { left: -48px; top: -3340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Cs2axe-vhhrIe { left: -40px; top: -2222px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-J6RZ7b { left: -62px; top: -1062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S { left: -40px; top: -3574px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S-r9oPif { left: 0px; top: -1912px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-IbE0S-i5vt6e { left: -40px; top: -1544px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-RWgCYc-yY4Wcc { left: -62px; top: -12938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-RWgCYc-yY4Wcc-BHsdwc { left: 0px; top: -6126px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-uiYelc { left: -40px; top: -10486px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NBDE7b-JaPV2b { left: -42px; top: -12668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-yHKmmc { left: 0px; top: -9472px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-yHKmmc-E3DyYd { left: -40px; top: -6872px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-hgHJW { left: 0px; top: -9300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-hgHJW-E3DyYd { left: -20px; top: -3996px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-lm6F6 { left: -22px; top: -2528px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-lm6F6-E3DyYd { left: 0px; top: -10716px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-X808Kb { left: -52px; top: -1872px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-X808Kb-E3DyYd { left: -22px; top: -4670px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-BvBYQ { left: 0px; top: -12526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-BvBYQ-E3DyYd { left: -42px; top: -5492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-tSZMSb { left: -40px; top: -2774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-An9n3c-tSZMSb-E3DyYd { left: 0px; top: -1718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q0hgme-mSEUvf { left: -40px; top: -5388px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-jyrRxf { left: 0px; top: -8454px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MHYjYb-nKQ6qf { left: 0px; top: -6896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RPzgNd-vfifzc-RxYbNe { left: 0px; top: -8650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-E8fGCc { left: 0px; top: -5988px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-t6UvL { left: -20px; top: -9300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-cGMI2b { left: -26px; top: -10202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-LK5yu { left: -52px; top: -6564px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-qwU8Me { left: 0px; top: -11224px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g7W7Ed-VtOx3e-ma6Yeb { left: -26px; top: -8412px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-tsZdxf-HLvlvd { left: -62px; top: -1718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-T3iPGc-r9oPif { left: -40px; top: -3142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-zf3vf { left: 0px; top: -12102px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-zf3vf-r9oPif { left: 0px; top: -2456px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Jz7rA { left: -56px; top: -6428px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Jz7rA-r9oPif { left: -26px; top: -7818px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LIMNJb { left: -26px; top: -4754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KsV2dd-HLvlvd { left: -40px; top: -13074px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-QIk5de-OWB6Me-EFlEBf { left: -40px; top: -76px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ntN8G { left: -40px; top: -2918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RCfa3e { left: -62px; top: -7552px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd-HLvlvd { left: -42px; top: -11384px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd { left: -42px; top: -11344px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-bBybbf { left: -60px; top: -5514px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf { left: 0px; top: -7490px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-Xhs9z { left: -20px; top: -9014px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qPaVXd-yHKmmc { left: -62px; top: -10112px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qPaVXd-yHKmmc-MFS4be-u2z5K { left: -22px; top: -12860px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-km6h5c { left: 0px; top: -7058px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-km6h5c-i5vt6e-r9oPif { left: -26px; top: -10156px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-n8nH7-jyrRxf { left: 0px; top: -3142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-n8nH7-jyrRxf { left: 0px; top: -6362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c-QUIbkc-HLvlvd-GoS4Be { left: 0px; top: -9340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-feLNVc { left: 0px; top: -4126px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-feLNVc-r9oPif { left: -40px; top: -274px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe { left: -20px; top: -12102px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic { left: -62px; top: -300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-drxrmf-DKlKme { left: -42px; top: -4020px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-drxrmf-BvBYQ { left: -22px; top: -1396px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ReqAjb-XaHFse { left: 0px; top: -12308px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb { left: -52px; top: -11104px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-E3Uge { left: -20px; top: -9034px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-ZdbLkb { left: -22px; top: -11000px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xceQUb-uPjwvb-ZdbLkb { left: 0px; top: -3340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g3I98d { left: -20px; top: -12840px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-elBQIf { left: -62px; top: -11694px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-vVewSc { left: -22px; top: -3842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-bMcfAe { left: -20px; top: -192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-oPu43-E3DyYd { left: -60px; top: -1478px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-oPu43-r9oPif { left: -26px; top: -9502px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-uDEFge-to915-r9oPif-oVleVe { left: -22px; top: -1370px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-i5vt6e-E3DyYd { left: -20px; top: -5492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-i5vt6e-r9oPif { left: 0px; top: -934px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e { left: -26px; top: -1934px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e-E3DyYd { left: -42px; top: -6654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-i5vt6e-r9oPif { left: 0px; top: -9420px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-i5vt6e-r9oPif { left: 0px; top: -8598px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-i5vt6e-E3DyYd { left: -20px; top: -8244px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-MFS4be-r9oPif-aOn1pf { left: 0px; top: -5044px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-i5vt6e-E3DyYd { left: -20px; top: -9206px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EnFNjd-i5vt6e-r9oPif { left: -22px; top: -13146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf-i5vt6e-E3DyYd { left: 0px; top: -2722px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-euCgFf-i5vt6e-r9oPif { left: 0px; top: -7032px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ihIZgd-i5vt6e-E3DyYd { left: 0px; top: -8324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HTJzpc-i5vt6e-E3DyYd { left: 0px; top: -4250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-w7bdYb { left: -26px; top: -8192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GEUYHe-r9oPif { left: -26px; top: -12328px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-r0zfL-HLvlvd { left: -42px; top: -10132px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe { left: -40px; top: -9972px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe { left: -20px; top: -212px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif { left: 0px; top: -7078px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif-v3pZbf { left: -34px; top: -9340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-r9oPif-HLvlvd { left: 0px; top: -8412px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P4Eybe-wcotoc-NkyfNe-uPjwvb-RvIlWb { left: -20px; top: -1084px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-CwllA-E3DyYd { left: 0px; top: -3280px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-E3Uge-E3DyYd { left: 0px; top: -13198px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-r9oPif { left: 0px; top: -4336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-HLvlvd-r9oPif { left: -26px; top: -5336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-r9oPif { left: -22px; top: -3340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-HLvlvd-r9oPif { left: -52px; top: -10202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-hgHJW-r9oPif { left: 0px; top: -582px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-yHKmmc-r9oPif { left: -46px; top: -1518px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-r9oPif { left: -48px; top: -7464px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc-E3Uge-r9oPif { left: 0px; top: -9854px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nEeMgc { left: -22px; top: -11284px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RFAvhb-jyrRxf-r9oPif { left: 0px; top: -4374px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-r9oPif { left: -20px; top: -11224px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-auswjd-r9oPif { left: -52px; top: -6606px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-Xhs9z-r9oPif { left: 0px; top: -252px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VPIWce-E3DyYd { left: 0px; top: -10978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ { left: -60px; top: -9380px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ-E3DyYd { left: 0px; top: -12668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JK9eJ-RvIlWb { left: -52px; top: -9092px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-ibnC6b { left: -20px; top: -8750px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XHoCPb-r9oPif-CwllA { left: -44px; top: -8832px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sfGayb-jbwjpc { left: 0px; top: -3512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-N7Eqid-W3lGp { left: -58px; top: -12250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-H8nU8b-W3lGp { left: -16px; top: -5004px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VgQDD-RPzgNd-vfifzc-RxYbNe-W3lGp { left: -26px; top: -7910px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rymPhb-r9oPif { left: -26px; top: -6696px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-kODWGd { left: 0px; top: -1172px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ndfHFb-yEEHq { left: 0px; top: -8670px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ge6pde-LkdAo-QG5zS { left: 0px; top: -8516px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pI3EI { left: -40px; top: -12360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e { left: -20px; top: -3040px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-nQ1Faf-E3DyYd { left: 0px; top: -5804px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-E3DyYd { left: 0px; top: -2896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-HLvlvd { left: -40px; top: -9992px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-nUpftc-YuD1xf { left: -20px; top: -300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-nUpftc-YuD1xf-IT5dJd-iBxYy-hxXJme-AHe6Kc { left: -22px; top: -6382px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf { left: -40px; top: -2938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf-IT5dJd-iBxYy-hxXJme-AHe6Kc { left: 0px; top: -12754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eMXQ4e-jNm5if-YuD1xf-mPlZac { left: -22px; top: -12668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc { left: 0px; top: -11738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc-HLvlvd { left: 0px; top: -8150px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-pGuBYc-FNFY6c { left: -22px; top: -4400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { left: 0px; top: -10506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY-r9oPif { left: 0px; top: -7672px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-p2N3pf-r9oPif { left: -22px; top: -12184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-N7Eqid { left: -22px; top: -4628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-DcLNVc-r9oPif { left: 0px; top: -9092px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-hgHJW { left: -34px; top: -5004px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-yHKmmc { left: -62px; top: -10268px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c-E3Uge { left: -52px; top: -11022px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ij8cu-E3Uge { left: -62px; top: -3594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc-uFfGwd { left: -52px; top: -6498px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JNdkSc { left: -42px; top: -6126px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-iMG1U-E3Uge { left: 0px; top: -12486px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GSQQnc-c4YZDc-r9oPif-HLvlvd { left: 0px; top: -6696px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ugYG9-c4YZDc { left: -20px; top: -11264px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ugYG9-c4YZDc-r9oPif-HLvlvd { left: 0px; top: -7646px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc-r9oPif-HLvlvd { left: -42px; top: -2528px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jCCvxc-r9oPif-HLvlvd { left: 0px; top: -7890px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk { left: -60px; top: -3574px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-rYk4U { left: 0px; top: -3492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-oScmOd { left: -20px; top: -4848px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-oScmOd { left: 0px; top: -12142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-oScmOd { left: 0px; top: -5216px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-FMvwCe-oScmOd { left: -20px; top: -320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-FMvwCe-oScmOd { left: 0px; top: -12938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-FMvwCe-oScmOd { left: 0px; top: -2180px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-HB1eCd-u2z5K { left: -22px; top: -9054px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-RFAvhb-u2z5K { left: -20px; top: -11900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-a1e4Ad-u2z5K { left: 0px; top: -6276px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-QymXn-u2z5K { left: -26px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-JeMQb { left: 0px; top: -10548px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-JeMQb { left: 0px; top: -1274px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-JeMQb { left: 0px; top: -2648px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-JeMQb { left: 0px; top: -12980px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-JeMQb { left: 0px; top: -7188px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-fmcmS { left: -40px; top: -608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-i8xkGf-fmcmS { left: -42px; top: -10290px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-fmcmS { left: -42px; top: -9634px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-LhcNjd-fmcmS { left: -20px; top: -5106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-SfQLQb-fmcmS { left: -60px; top: -7012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-TzA9Ye-SfQLQb-fmcmS { left: -22px; top: -3452px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-fmcmS { left: -52px; top: -6632px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-KLRBe-fmcmS { left: -40px; top: -1658px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-fmcmS { left: -22px; top: -12002px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .VIpgJd-INgbqf-LgbsSe-barxie .HB1eCd-Bz112c-fmcmS-efjR6d-gNy6Jf-fmcmS { left: 0px; top: -5258px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-LK5yu-Ysl7Fe { left: 0px; top: -8350px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-oXtfBe-Ysl7Fe { left: 0px; top: -4566px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-ma6Yeb-qwU8Me-Ysl7Fe { left: 0px; top: -11592px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-LK5yu-Ysl7Fe { left: -26px; top: -952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-Ysl7Fe { left: 0px; top: -8878px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-oXtfBe-qwU8Me-Ysl7Fe { left: 0px; top: -5408px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-LK5yu-Ysl7Fe { left: -26px; top: -4500px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-oXtfBe-Ysl7Fe { left: 0px; top: -11048px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-mAKE4e-neVct-cGMI2b-qwU8Me-Ysl7Fe { left: -26px; top: -11428px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qknJed-AFZkUd { left: 0px; top: -4060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-qknJed-AFZkUd-hJDwNd { left: -62px; top: -3642px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JLm1tf-DJPBic-AFZkUd-W3lGp-TLxrU { left: -46px; top: -3804px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RFnRab-r9oPif { left: 0px; top: -10690px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd { left: -60px; top: -3040px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc { left: -42px; top: -3452px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-aOn1pf { left: -20px; top: -4272px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-VqDHhd { left: -62px; top: -10092px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc { left: -62px; top: -1150px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc-E3DyYd { left: -20px; top: -3080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me { left: -20px; top: -6722px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-aOn1pf { left: -20px; top: -7146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd-r9oPif { left: -48px; top: -1892px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-r9oPif { left: 0px; top: -2998px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-di8rgd-aSWTkc-r9oPif-aOn1pf { left: 0px; top: -2502px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-r9oPif-VqDHhd { left: -52px; top: -4080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Vj7tjb-SYBOGc-r9oPif { left: -22px; top: -13094px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-r9oPif { left: -46px; top: -11124px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-OWB6Me-r9oPif-aOn1pf { left: 0px; top: -556px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb { left: 0px; top: -2072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-JaPV2b { left: 0px; top: -960px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-r9oPif { left: -55px; top: -5086px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XHgP6b-dNswIb-r9oPif-gS7Ybc { left: 0px; top: -6830px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG { left: 0px; top: -9280px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-r9oPif { left: -52px; top: -1846px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-MFS4be-ETmUib { left: 0px; top: -5470px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-SeBwEf { left: -26px; top: -7844px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-SeBwEf-r9oPif { left: -20px; top: -4166px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b { left: -20px; top: -1478px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-GjlSrc { left: 0px; top: -648px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-V7AMae { left: -20px; top: -12820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-CwllA { left: 0px; top: -1544px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ONu0F { left: 0px; top: -8556px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-r9oPif { left: 0px; top: -2800px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-i5vt6e-TY4T7c { left: -20px; top: -4650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-E3DyYd { left: -20px; top: -12572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-r9oPif { left: -26px; top: -12728px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-r9oPif { left: -22px; top: -3616px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d { left: -42px; top: -6456px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-r9oPif { left: 0px; top: -882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq { left: -62px; top: -7532px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-VtOx3e { left: 0px; top: -1678px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-MFS4be { left: 0px; top: -76px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-Q4BLdf { left: -20px; top: -8476px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-r9oPif { left: 0px; top: -10012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hSRGPd-di8rgd-r9oPif { left: -42px; top: -3202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-Hjleke-r9oPif { left: 0px; top: -5336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ft5J4b-iOyk4d-r9oPif { left: 0px; top: -4520px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-bVEB4e { left: -20px; top: -12230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nGOfy-Dy7EIf { left: -52px; top: -2046px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YRhSCb-Dy7EIf { left: -42px; top: -3996px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ryxqyc-vUjI9d-hxGuWb { left: 0px; top: -484px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ryxqyc-pDPzzb-hxGuWb { left: -40px; top: -5086px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-muPwQb { left: -35px; top: -484px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-x5cW0b { left: 0px; top: -11778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-ma6Yeb-LK5yu { left: 0px; top: -5926px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-cXXICe-ma6Yeb-qwU8Me { left: 0px; top: -3452px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-vbnc8b { left: 0px; top: -4106px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-vbnc8b-r9oPif { left: -52px; top: -9538px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-r9oPif { left: -20px; top: -9228px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-r9oPif-HLvlvd { left: 0px; top: -9906px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-Qs3R8d-RvIlWb { left: -52px; top: -556px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-Qs3R8d-RvIlWb { left: -40px; top: -5608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-uPjwvb-RvIlWb { left: -52px; top: -9808px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-uPjwvb-RvIlWb { left: 0px; top: -12546px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-r9oPif { left: 0px; top: -10156px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-LSK72c-r9oPif { left: -26px; top: -7378px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-jNm5if-LrF0Pc-r9oPif { left: 0px; top: -4080px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-r9oPif { left: -26px; top: -8594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-tcqZEf-r9oPif { left: -46px; top: -7844px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DfC5c-UVuwbd-LrF0Pc-r9oPif { left: 0px; top: -2376px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YxWbQd-r9oPif { left: 0px; top: -908px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YxWbQd { left: -20px; top: -3320px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb { left: 0px; top: -4650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-ZdbLkb { left: 0px; top: -10896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-uPjwvb-ZdbLkb { left: 0px; top: -7464px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-QLEXN-ZdbLkb { left: -52px; top: -7820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-wvGCSb-LoDsGd-jJ3Q2c-Q7Syqe-r9oPif { left: 0px; top: -11428px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jEEo8-HLvlvd { left: -20px; top: -8130px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RxTQ8e-oq6NAc { left: -26px; top: -4374px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Y5dbrb-r9oPif { left: -26px; top: -12546px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KNM5Ef { left: -40px; top: -3684px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue { left: -26px; top: -5044px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue-r9oPif { left: 0px; top: -9254px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-H6hmue-RAze1d-r9oPif { left: -22px; top: -7464px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-r9oPif-aOn1pf { left: 0px; top: -7398px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-clhnwb { left: -40px; top: -8536px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e4raY { left: 0px; top: -9952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-rYk4U { left: -40px; top: -7012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vOBb1e { left: -40px; top: -2436px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-smkJ3e { left: 0px; top: -12360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YJL97b { left: -62px; top: -4250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YJL97b-r9oPif { left: -46px; top: -8192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-tSZMSb { left: -40px; top: -9952px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-m3mY0d-RbRzK { left: -44px; top: -9696px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PZMiD-M1QMZb-fmcmS { left: -20px; top: -10958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YLEF4c { left: -20px; top: -4146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb { left: -58px; top: -170px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-W3lGp { left: 0px; top: -6762px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-E3DyYd { left: -40px; top: -5874px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-F9IAbd-HSrbLb-r9oPif { left: -46px; top: -12400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-Wz3zdc-Z7HxEc-r9oPif-T60B1 { left: -26px; top: -8218px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-Wz3zdc-Z7HxEc-LrF0Pc-r9oPif { left: 0px; top: -5186px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-hWJfub-yHKmmc-r9oPif-T60B1 { left: -26px; top: -9118px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-oSWire { left: -40px; top: -5470px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe { left: -22px; top: -4250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-E3DyYd { left: -22px; top: -9696px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-r9oPif { left: -22px; top: -13172px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-z5C9Gb-P5Aqpe-Qs3R8d-RvIlWb { left: 0px; top: -10202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Faem2b-cVFi4-r9oPif-mPlZac { left: 0px; top: -5362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-V67aGc-i5vt6e { left: 0px; top: -6028px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-MPu53c-C2S4ob { left: 0px; top: -2114px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd-G0jgYd-r9oPif { left: 0px; top: -6250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-n6j7Re { left: -40px; top: -232px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uaxL4e-n6j7Re { left: 0px; top: -1478px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-h976Ve { left: -46px; top: -7646px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-ctOWCc-r9oPif { left: -48px; top: -9420px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eizL8e-Vgu1H-r9oPif { left: -26px; top: -2154px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-npMLoc-r9oPif { left: -20px; top: -11124px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop { left: 0px; top: -4272px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-E3DyYd { left: 0px; top: -4314px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-r9oPif { left: -46px; top: -10622px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-SIsrTd { left: -20px; top: -6048px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Gbxop-SIsrTd-E3DyYd { left: 0px; top: -8812px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe { left: 0px; top: -9654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-HLvlvd { left: -26px; top: -4314px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-zYyPae { left: 0px; top: -13136px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-GjlSrc { left: 0px; top: -2222px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-V7AMae { left: -20px; top: -7424px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-uQPRwe-CwllA { left: -42px; top: -11324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-gNuiOc-r9oPif { left: -26px; top: -9092px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-gNuiOc-HLvlvd-r9oPif { left: -46px; top: -836px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed { left: -20px; top: -2094px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-lQVAed-r9oPif { left: 0px; top: -7598px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-clPPge-r9oPif { left: -26px; top: -5900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-clPPge-E3DyYd { left: -40px; top: -3594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-r9oPif { left: -48px; top: -13142px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-u5Azmc { left: -20px; top: -6362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-LBRlSe { left: 0px; top: -12440px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GnPzId { left: -20px; top: -232px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-xZDoyc-MJ0UK { left: -40px; top: -12506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-a2ItGd { left: 0px; top: -13054px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-wWDucd { left: -40px; top: -4650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GEUYHe { left: -20px; top: -7012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-WX1Rmf { left: -20px; top: -3060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-c6tfMc { left: 0px; top: -3554px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e3uGsb { left: -40px; top: -2114px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-e3uGsb-C2NXRc { left: -40px; top: -10446px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VkLyEc { left: -26px; top: -9854px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-I3TTMc { left: -60px; top: -9340px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-I3TTMc-nQ1Faf { left: -20px; top: -1658px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-r9oPif { left: -52px; top: -10922px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-E3DyYd { left: -20px; top: -5708px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-nUpftc-mG3Az-r9oPif { left: -52px; top: -11618px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-bstyQc { left: -20px; top: -2938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-u5Azmc-r9oPif { left: 0px; top: -9512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-LBRlSe-r9oPif { left: -52px; top: -12774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GnPzId-r9oPif { left: 0px; top: -11022px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-xZDoyc-MJ0UK-r9oPif { left: 0px; top: -8192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-a2ItGd-r9oPif { left: -22px; top: -1820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-wWDucd-r9oPif { left: 0px; top: -3228px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-GEUYHe-r9oPif { left: -52px; top: -10870px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-WX1Rmf-r9oPif { left: -46px; top: -8624px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wz3zdc-c6tfMc-r9oPif { left: -48px; top: -13116px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-hauLI-ETmUib { left: 0px; top: -11490px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-hauLI-r9oPif-ETmUib { left: -46px; top: -7672px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JEruSd-ETmUib { left: 0px; top: -5492px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-i4ewOd-r9oPif { left: -42px; top: -8324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-JEruSd-r9oPif-ETmUib { left: 0px; top: -9972px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-r9oPif { left: 0px; top: -8078px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-E3DyYd { left: 0px; top: -11654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H-uPjwvb-E3DyYd { left: -42px; top: -1778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-MFS4be-E3DyYd-t24pnf { left: 0px; top: -13094px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic-mlKF6d-kRWtF { left: 0px; top: -10052px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-J652Ic-LkdAo { left: -22px; top: -8324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-YjoMNe { left: -34px; top: -5968px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YjoMNe-IFdKyd { left: -20px; top: -842px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-YjoMNe-HLvlvd { left: 0px; top: -3882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-V5oUn { left: -20px; top: -8692px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vRvVU-wcotoc-xvr5H { left: -26px; top: -2416px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-h976Ve-r9oPif { left: -48px; top: -530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-YjoMNe-IFdKyd-r9oPif { left: -35px; top: -504px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-j4gsHd-hFsbo-bEDTcc-h976Ve { left: 0px; top: -1252px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-muPwQb-LSK72c-r9oPif { left: 0px; top: -8572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-iyXyEd { left: -48px; top: -5362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-LkdAo { left: 0px; top: -4500px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-u3p8pb-mzNpsf { left: 0px; top: -10622px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-iBxYy-Pv6Am { left: 0px; top: -4862px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jNm5if-DyVDA-r9oPif { left: -26px; top: -4774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-dZssN-D5MPn { left: 0px; top: -4780px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-g6cJHd-LkdAo-mPlZac { left: 0px; top: -2550px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-oSWire-r9oPif { left: 0px; top: -6606px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HB1eCd-F9IAbd-OVkoRd-yaNpec { left: -20px; top: -2134px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-r9oPif { left: -26px; top: -2046px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-r9oPif-HLvlvd { left: -48px; top: -3616px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-uPjwvb-RvIlWb { left: -52px; top: -12526px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-B8pEb-HLvlvd { left: -40px; top: -12082px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-zMQiGf-WAutxc { left: -40px; top: -10506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-SeDgR-V7AMae { left: -62px; top: -11364px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-t5jYtc-appOce { left: -46px; top: -4374px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TdyTDe-V7AMae { left: -26px; top: -12308px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DUGJie-appOce { left: 0px; top: -4984px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-aIWppb-htvI8d-r9oPif { left: -52px; top: -6538px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c { left: -40px; top: -2242px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-bOjP2c-u014N-ImhxVb-aTv5jf { left: -42px; top: -10112px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop { left: 0px; top: -688px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-SIsrTd { left: 0px; top: -436px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-B1neQd-i2RYZ { left: 0px; top: -10778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-ixlDHd-Gbxop-B1neQd-i2RYZ-SIsrTd { left: 0px; top: -6782px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nupQLb-J42Xof-zVpoTe { left: -40px; top: -1478px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-TIHSC-r9oPif { left: 0px; top: -2402px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TDvtud { left: -20px; top: -6856px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q3tln-x9Ufpf-SjW3R { left: -14px; top: -5926px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-rymPhb-Jn51gd-r9oPif { left: 0px; top: -4754px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-wcotoc-ndfHFb-E3DyYd { left: 0px; top: -1040px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DcLNVc-g6cJHd-E3DyYd { left: -42px; top: -794px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-ZdbLkb { left: -52px; top: -7798px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yEEHq-x5cW0b-E3DyYd { left: 0px; top: -12860px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Tswv1b-E3DyYd { left: 0px; top: -10334px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-VtOx3e-E3DyYd { left: -22px; top: -10978px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fI6EEc-MFS4be-E3DyYd-LSK72c { left: -61px; top: -504px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-DcLNVc-Xhs9z-E3DyYd { left: -42px; top: -5216px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-wUN2c-E3DyYd { left: 0px; top: -794px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-IAXTZb-E3DyYd { left: 0px; top: -9374px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Yygnk-E3DyYd { left: 0px; top: -2896px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Yygnk-Z5I80b-E3DyYd { left: -20px; top: -6654px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PrY1nf-UlP5cd-E3DyYd { left: -26px; top: -8572px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HB1eCd-DJPBic { left: 0px; top: -10738px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-a1e4Ad-DJPBic { left: 0px; top: -1396px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RFAvhb-DJPBic { left: -60px; top: -12360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Poonxc-eEGnhe { left: -20px; top: -1678px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Poonxc-eEGnhe-r9oPif { left: -52px; top: -4796px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nyE0bc-r9oPif { left: -46px; top: -2482px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-E3DyYd { left: -58px; top: -11900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-LK5yu-E3DyYd { left: -22px; top: -10736px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-qwU8Me-E3DyYd { left: -42px; top: -7104px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Q8Kwad-hgHJW-E3DyYd { left: -26px; top: -9420px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-OCFbXc-E3DyYd { left: 0px; top: -9694px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-z5C9Gb-E3DyYd { left: -52px; top: -10848px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xl07Ob-E3DyYd { left: -20px; top: -7512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WAutxc-jNm5if-MFS4be-E3DyYd { left: -46px; top: -4334px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-OiiCO-E3DyYd { left: 0px; top: -8104px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-nUpftc-E3DyYd { left: 0px; top: -4800px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ObfsIf-nUpftc-MFS4be-E3DyYd { left: -40px; top: -11694px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-u0pjoe-MFS4be-ETmUib { left: 0px; top: -2918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-E3DyYd { left: -26px; top: -5362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-KqJenf-nllRtd-E3DyYd { left: -38px; top: -6276px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-uPjwvb-ZdbLkb { left: -26px; top: -7772px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-j4gsHd-IT5dJd-XxIAqe-E3DyYd { left: 0px; top: -3202px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-E3DyYd { left: -20px; top: -10668px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-xAa0Lb-ShBeI-E3DyYd { left: -40px; top: -5660px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Fs2VSc-r9oPif { left: 0px; top: -7772px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TNZ3Zd { left: -62px; top: -11838px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TNZ3Zd-r9oPif { left: -52px; top: -582px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-yaNpec { left: 0px; top: -1698px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TZk80d-jCCvxc-HNJgkc { left: -60px; top: -4650px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Bpn8Yb-E3DyYd { left: 0px; top: -11324px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-aTv5jf-km6h5c-jirZld-r9oPif { left: 0px; top: -6520px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-UlP5cd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HivRGb-ZlOZYc-UlP5cd { left: 0px; top: -11550px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-JbbQac-E3DyYd { left: -22px; top: -7490px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-kWbB0e-kWTbQe-E3DyYd { left: -46px; top: -3778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-n5AaSd-E3DyYd { left: -52px; top: -10730px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rsbfue-E3DyYd { left: -46px; top: -9232px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-VtOx3e-hxXJme-E3DyYd { left: 0px; top: -1230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ayzxhb-XPtOyb-r9oPif { left: -26px; top: -11022px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-PLDbbf-Ysl7Fe-XZYQce { left: 0px; top: -10356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-PLDbbf-SIsrTd-Ysl7Fe-XZYQce { left: 0px; top: -3382px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-DARUcf-n5AaSd-Ysl7Fe-XZYQce { left: -22px; top: -5804px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-DARUcf-n5AaSd-SIsrTd-Ysl7Fe-XZYQce { left: -26px; top: -5146px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hFsbo-NGme3c-yY4Wcc-E3DyYd { left: 0px; top: -8770px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-eEDwDf-xSh02c-E3DyYd { left: 0px; top: -11000px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XPtOyb-VFQeR-E3DyYd { left: -22px; top: -8812px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-kWbB0e-kWTbQe-E3DyYd { left: 0px; top: -1778px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-ltEGzf-E3DyYd { left: 0px; top: -12022px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-RPzgNd-E3DyYd { left: 0px; top: -9446px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Wxxdob-fmcmS-i8xkGf-E3DyYd { left: 0px; top: -7624px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Ge5tnd-fmcmS-E3DyYd { left: -58px; top: -2570px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-E3DyYd { left: 0px; top: -3616px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-E3DyYd { left: -26px; top: -6540px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-MFS4be-E3DyYd { left: -42px; top: -3512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-hFsbo-FMODoe-E3DyYd { left: -46px; top: -10012px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-LkdAo-E3DyYd { left: 0px; top: -1820px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-LkdAo-MFS4be-E3DyYd { left: -48px; top: -12162px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-dajHKf-E3DyYd { left: 0px; top: -4442px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-dajHKf-MFS4be-E3DyYd { left: -52px; top: -10826px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-BaYisc-E3DyYd { left: -26px; top: -9880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-CpWD9d-BaYisc-MFS4be-E3DyYd { left: -60px; top: -1438px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-E3DyYd { left: -44px; top: -9586px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-E3DyYd { left: -20px; top: -10290px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-MFS4be-E3DyYd { left: -40px; top: -6742px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-hFsbo-FMODoe-E3DyYd { left: 0px; top: -1416px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-LkdAo-E3DyYd { left: -22px; top: -1348px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-LkdAo-MFS4be-E3DyYd { left: -60px; top: -1544px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-dajHKf-E3DyYd { left: -60px; top: -9184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-dajHKf-MFS4be-E3DyYd { left: 0px; top: -9586px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-BaYisc-E3DyYd { left: -44px; top: -11000px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-RWgCYc-I3Yihd-BaYisc-MFS4be-E3DyYd { left: 0px; top: -12184px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TDvtud-r9oPif { left: -22px; top: -9608px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-G0jgYd-E3DyYd-EnQdTb { left: -26px; top: -7078px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-hPL1Ee-Ysl7Fe-XZYQce { left: -26px; top: -882px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Rgqkje-hPL1Ee-SIsrTd-Ysl7Fe-XZYQce { left: 0px; top: -10826px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-LK5yu-JeMQb { left: 0px; top: -12594px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-oXtfBe-JeMQb { left: 0px; top: -7262px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-qwU8Me-JeMQb { left: 0px; top: -11150px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-LK5yu-JeMQb { left: 0px; top: -1958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-JeMQb { left: 0px; top: -5730px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-qwU8Me-JeMQb { left: 0px; top: -8940px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-LK5yu-JeMQb { left: 0px; top: -2262px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-oXtfBe-JeMQb { left: 0px; top: -96px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-qwU8Me-JeMQb { left: 0px; top: -362px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-LK5yu-t5QKTe { left: 0px; top: -8266px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-oXtfBe-t5QKTe { left: 0px; top: -2570px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-ma6Yeb-qwU8Me-t5QKTe { left: 0px; top: -5278px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-LK5yu-t5QKTe { left: 0px; top: -736px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-t5QKTe { left: 0px; top: -6068px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-oXtfBe-qwU8Me-t5QKTe { left: 0px; top: -12250px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-LK5yu-t5QKTe { left: 0px; top: -4192px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-oXtfBe-t5QKTe { left: -22px; top: -4442px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-mAKE4e-neVct-cGMI2b-qwU8Me-t5QKTe { left: -20px; top: -1172px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-LK5yu-KW5YQd-JeMQb { left: 0px; top: -6938px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-oXtfBe-KW5YQd-JeMQb { left: 0px; top: -1584px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-qwU8Me-KW5YQd-JeMQb { left: 0px; top: -3922px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-efjR6d-TzA9Ye-JeMQb { left: 0px; top: -7930px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-efjR6d-i8xkGf-JeMQb { left: 0px; top: -7698px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-aP0wEc-JeMQb { left: 0px; top: -8004px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-LK5yu-JeMQb { left: 0px; top: -5534px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-jyrRxf-fmcmS-i8xkGf-mhHukc-qwU8Me-JeMQb { left: 0px; top: -3704px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-s2ctBd-E3DyYd { left: -26px; top: -530px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-r9oPif { left: 0px; top: -8624px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-w9NWI-r9oPif { left: -26px; top: -10690px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-z5C9Gb { left: 0px; top: -5708px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-OCFbXc { left: 0px; top: -3996px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-tJHJj { left: -60px; top: -76px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-tJHJj-r9oPif { left: -40px; top: -9014px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-tJHJj { left: -20px; top: -7356px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-tJHJj-r9oPif { left: -52px; top: -7378px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-vhaaFf-J9pn5c-r9oPif { left: 0px; top: -5874px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-KoToPc-J9pn5c-r9oPif { left: 0px; top: -12774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd-E3DyYd { left: -40px; top: -6850px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-yOOK0-IFdKyd-MFS4be-E3DyYd { left: -22px; top: -9586px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-l4eHX-t0O9Gd-XpSwdc { left: -42px; top: -1130px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-EWK8Bb-lxyxlb-XpSwdc { left: 0px; top: -10228px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-MFS4be-ZdbLkb { left: -52px; top: -11062px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-MFS4be-uPjwvb-ZdbLkb { left: -26px; top: -1912px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GhbEaf-xFQqWe-RvIlWb { left: -52px; top: -3228px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-ZdbLkb { left: -34px; top: -5946px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-uPjwvb-ZdbLkb { left: 0px; top: -4628px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-RvIlWb { left: 0px; top: -10072px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-WSzvjf-uPjwvb-RvIlWb { left: 0px; top: -6336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-yqoORe-XpSwdc { left: -20px; top: -12082px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HrRdod-yLHjwb-yqoORe-RvIlWb { left: -20px; top: -4890px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-Jw1b8-uPjwvb-r9oPif { left: -22px; top: -8104px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-XPtOyb-VFQeR-XpSwdc { left: -20px; top: -2918px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-pGuBYc-ZdbLkb { left: -20px; top: -8454px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PGTmtf-ZdbLkb { left: 0px; top: -1370px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nLfZJb-r9oPif { left: 0px; top: -9880px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fcEm8e-r9oPif { left: -56px; top: -5926px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-CSqGDb-yaNpec { left: 0px; top: -2336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-E3DyYd { left: -60px; top: -4292px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-flHhI-fmcmS-CSqGDb-r9oPif { left: -26px; top: -12774px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nctj2d-yaNpec { left: -26px; top: -2376px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nctj2d-E3DyYd { left: -60px; top: -2222px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-g5XWbe-yaNpec { left: -20px; top: -8712px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HiaYvf-g5XWbe-r9oPif { left: 0px; top: -7818px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-sA2X9e-KbLeYb-E3DyYd { left: -26px; top: -1034px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LUSEYe { left: 0px; top: -11900px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-LUSEYe-J9pn5c-r9oPif { left: 0px; top: -2154px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-h1U9Be { left: -62px; top: -12958px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DyVDA-h1U9Be-J9pn5c-r9oPif { left: -20px; top: -816px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-HLvlvd-r9oPif { left: -22px; top: -9718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-HLvlvd-r9oPif { left: -52px; top: -9512px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-HLvlvd-i5vt6e-r9oPif { left: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-HLvlvd-i5vt6e-r9oPif { left: -26px; top: -9828px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-mrxPge-r9oPif { left: 0px; top: -3254px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-mrxPge-r9oPif { left: 0px; top: -12334px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-yHKmmc-mrxPge-i5vt6e-r9oPif { left: 0px; top: -1846px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-hWJfub-hgHJW-mrxPge-i5vt6e-r9oPif { left: -22px; top: -9446px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-h9d3hd-E3DyYd { left: -48px; top: -1396px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-Vkfede-ZdbLkb { left: 0px; top: -3466px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-TvD9Pc-n9oEIb-ZdbLkb { left: 0px; top: -9718px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P8wAXc-wcotoc-XzMRXd-XpSwdc { left: -52px; top: -8898px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-P8wAXc-wcotoc-XzMRXd-RvIlWb { left: 0px; top: -1518px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-FNFY6c-bEDTcc-HzdVzc-RvIlWb { left: 0px; top: -12728px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-hFsbo-XpSwdc { left: -42px; top: -3280px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-NziyQe-hFsbo-HLvlvd-XpSwdc { left: -20px; top: -12506px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HvfI2b-XpSwdc { left: -42px; top: -3862px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-HvfI2b-HLvlvd-XpSwdc { left: -22px; top: -794px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-uPjwvb-ZdbLkb { left: -22px; top: -11838px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-htvI8d-uPjwvb-RvIlWb { left: -52px; top: -6336px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-RvIlWb { left: -26px; top: -1846px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-ZdbLkb { left: 0px; top: -11716px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-fQQGY-XpSwdc { left: 0px; top: -12230px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c-E3DyYd { left: 0px; top: -4400px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-nKQ6qf-Y80K8c-r9oPif { left: 0px; top: -10446px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-GMvhG-FFXbQc-ZdbLkb { left: -26px; top: -8432px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-yHKmmc-XpSwdc { left: 0px; top: -8536px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-PFprWc-hgHJW-XpSwdc { left: -40px; top: -4060px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ImhxVb-nMj4jb-xFQqWe-ZdbLkb { left: 0px; top: -278px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-ImhxVb-nMj4jb-MFS4be-ZdbLkb { left: -52px; top: -6584px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c-DJPBic-v3pZbf-ZdbLkb { left: -20px; top: -4020px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c { direction: ltr; text-align: left; height: 60px; overflow: hidden; vertical-align: middle; width: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/branding_sprite1.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-RJLb9c { position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-ndfHFb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-zTETae { left: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-TftRv { left: 0px; top: -180px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-G1jlMc { left: 0px; top: -300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-arrpzb { left: 0px; top: -360px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-QymXn { left: 0px; top: -60px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-t02dhe { left: 0px; top: -120px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-n7vHCb-Bz112c-jdTLZc { left: 0px; top: -240px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c { direction: ltr; text-align: left; height: 21px; overflow: hidden; vertical-align: middle; width: 21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/jfk_sprite186.png"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-RJLb9c-VVu2ae { }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c-RJLb9c-haAclf { height: 4167px; position: absolute; width: 42px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-hxXJme-xl07Ob-LgbsSe-uDEFge .HB1eCd-Bz112c { height: 19px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-RJLb9c-haAclf { opacity: 0.55; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-OMz1o, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-usbjsf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-EgTfg, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-hDEnYe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-I9GLp, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-nA1mMd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-wlNA0d, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c .HB1eCd-Bz112c-jSFuyb { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-jCCvxc-hSRGPd { width: 500px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .jCCvxc-hSRGPd-Sx9Kwc { color: black; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; white-space: normal; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .jCCvxc-hSRGPd-PLEiK-ZYyEqf { position: absolute; top: 0px; padding-top: 16px; left: 220px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble { border: 1px solid rgb(238, 238, 238); box-shadow: rgba(0, 0, 0, 0.05) 0px 3px 3px; background: rgba(255, 255, 255, 0.85); border-radius: 41px; position: absolute; top: 0px; width: 40px; text-align: center; z-index: -2; cursor: default; opacity: 0; transition: opacity 0.25s ease-in-out 0s, z-index 0.26s linear 0.25s; transform: translate(-50%, -50%); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble.RXQi4b-tiLKmf-RCfa3e { z-index: 101; visibility: hidden; transition: visibility 0s linear 0.25s, opacity 0.25s ease-in-out 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble.HB1eCd-DfC5c-VCkuzd-ZiwkRe { opacity: 1; cursor: pointer; z-index: 101; transition: opacity 0.25s ease-in-out 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble.HB1eCd-DfC5c-VCkuzd-ZiwkRe.RXQi4b-tiLKmf-RCfa3e { visibility: visible; transition-delay: 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble.HB1eCd-DfC5c-VCkuzd-mAKE4e-ZYIfFd { z-index: -2; opacity: 0; top: 0px; transition: none 0s ease 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble.HB1eCd-DfC5c-VCkuzd-mAKE4e-ZYIfFd.RXQi4b-tiLKmf-RCfa3e { z-index: 101; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble:hover { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble:focus { outline: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble .HB1eCd-DfC5c-VCkuzd-haAclf { border-radius: 41px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble .DfC5c-LgbsSe.r08add-ZiwkRe-LgbsSe { border-top-left-radius: 41px; border-top-right-radius: 41px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-instant-bubble .DfC5c-LgbsSe.E6eRQd-ZiwkRe-LgbsSe { border-bottom-left-radius: 41px; border-bottom-right-radius: 41px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf #docs-instant-bubble { background: rgb(249, 251, 253); border: none; box-shadow: rgba(0, 0, 0, 0.15) 0px 4px 8px 3px, rgba(0, 0, 0, 0.3) 0px 1px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .DPvwYc { font-family: "Material Icons Extended"; font-weight: normal; font-style: normal; font-size: 24px; line-height: 1; letter-spacing: normal; text-rendering: optimizelegibility; text-transform: none; display: inline-block; overflow-wrap: normal; direction: ltr; font-feature-settings: "liga"; -webkit-font-smoothing: antialiased; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb html[dir="rtl"] .sm8sCf { transform: scaleX(-1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c { border: 2px solid rgb(95, 99, 104); border-radius: 2px; box-sizing: border-box; cursor: pointer; height: 18px; margin: 1px; outline: none; flex-shrink: 0; top: 4px; width: 18px; display: inline-block; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd { background-color: rgb(26, 115, 232); border: 2px solid rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iI2ZmZiIvPjwvc3ZnPg=="); display: block; line-height: 15px; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iQ2FudmFzVGV4dCIvPjwvc3ZnPg=="); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd::before { border-top: 2px solid white; content: ""; display: block; height: 0px; margin-left: 3px; margin-top: 6px; width: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { border: 2px solid rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me { cursor: default; opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie { background-clip: padding-box; background-color: rgb(95, 99, 104); border-color: rgb(95, 99, 104); opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { background-color: rgb(26, 115, 232); border: 2px solid rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-uE9yNd { background-clip: padding-box; background-color: rgb(95, 99, 104); border-color: rgb(95, 99, 104); opacity: 0.38; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-MPu53c-LkdAo, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-MPu53c-LkdAo { background-color: highlight; opacity: 0.38; z-index: -1; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb span.HB1eCd-HzV7m-UMrnmb-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie { border-color: graytext; opacity: 1; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c { -webkit-box-align: start; align-items: flex-start; cursor: pointer; display: flex; max-width: 672px; outline: none; padding: 8px 0px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-bN97Pc { flex-shrink: 1; margin-left: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { width: 40px; height: 40px; border-radius: 50%; cursor: pointer; margin-left: -10px; margin-top: -10px; position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c { border: 2px solid rgb(95, 99, 104); border-radius: 2px; box-sizing: border-box; cursor: pointer; height: 18px; margin: 1px; outline: none; flex-shrink: 0; top: 4px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-uE9yNd { background-color: rgb(26, 115, 232); border: 2px solid rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iI2ZmZiIvPjwvc3ZnPg=="); display: block; line-height: 15px; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iQ2FudmFzVGV4dCIvPjwvc3ZnPg=="); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-uE9yNd::before { border-top: 2px solid white; content: ""; display: block; height: 0px; margin-left: 3px; margin-top: 6px; width: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c { cursor: default; opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ZmdkE .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.04; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.06; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-uE9yNd { background-clip: padding-box; background-color: rgb(95, 99, 104); border-color: rgb(95, 99, 104); opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ZmdkE .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie + .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.04; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie + .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.06; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie + .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-V67aGc { color: rgb(60, 64, 67); cursor: pointer; display: block; font: 14px / 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 3px 0px; width: auto; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-V67aGc { cursor: default; opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ij8cu { color: rgb(95, 99, 104); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; padding: 1px 0px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ij8cu { opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ij8cu-ZYIfFd { display: none; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie + .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie + .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-LkdAo { background-color: highlight; opacity: 0.38; z-index: -1; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-barxie { border-color: graytext; opacity: 1; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-V67aGc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c.HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-xO8zKb-MPu53c-ij8cu { color: graytext; opacity: 1; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c { -webkit-box-align: start; align-items: flex-start; cursor: pointer; display: flex; max-width: 672px; outline: none; padding: 8px 0px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { width: 40px; height: 40px; border-radius: 50%; cursor: pointer; margin-left: -10px; margin-top: -10px; position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c { border: 2px solid rgb(95, 99, 104); border-radius: 2px; box-sizing: border-box; cursor: pointer; height: 18px; margin: 1px; outline: none; flex-shrink: 0; top: 4px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-uE9yNd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c { background-color: rgb(26, 115, 232); border: 2px solid rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iI2ZmZiIvPjwvc3ZnPg=="); display: block; line-height: 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-uE9yNd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c::before { border-top: 2px solid white; content: ""; display: block; height: 0px; margin-left: 3px; margin-top: 6px; width: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c { cursor: default; opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-ZmdkE .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.04; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.06; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(95, 99, 104); opacity: 0.1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-uE9yNd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c { background-clip: padding-box; background-color: rgb(95, 99, 104); border-color: rgb(95, 99, 104); opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-ZmdkE.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.04; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-XpnDCe.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.06; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-auswjd.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: rgb(26, 115, 232); opacity: 0.1; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c::before { content: url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHZpZXdCb3g9IjAgMCAxIDEiIHByZXNlcnZlQXNwZWN0UmF0aW89InhNaW5ZTWluIG1lZXQiPjxwYXRoIGQ9Ik0uMDQuNjI3LjE0Ni41Mi40My44MDQuMzIzLjkxem0uMTc3LjE3N0wuODU0LjE2Ny45Ni4yNzMuMzIzLjkxeiIgZmlsbD0iQ2FudmFzVGV4dCIvPjwvc3ZnPg=="); }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-XpnDCe .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-auswjd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-LkdAo { background-color: highlight; opacity: 0.38; z-index: -1; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-barxie .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-OWB6Me.HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-uE9yNd .HB1eCd-HzV7m-UMrnmb-trycPc-MPu53c-MPu53c { border-color: graytext; opacity: 1; }
}

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { background: rgb(255, 255, 255); border: 1px solid transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; position: absolute; z-index: 1003; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); left: 0px; position: absolute; top: 0px; z-index: 998; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc:focus.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke { border-bottom: none; padding: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-fmcmS { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 22px; font-weight: 400; line-height: 28px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { height: 24px; position: absolute; right: 24px; top: 26px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-bN97Pc { min-width: 312px; padding: 0px 24px 24px; color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-c6xFrd { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 24px; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe, .HB1eCd-HzV7m-UMrnmb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe { text-transform: none; }

.HB1eCd-HzV7m-UMrnmb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-F75qrd-wcotoc-JIbuQc-LgbsSe.HB1eCd-HzV7m-LgbsSe { margin-left: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe { box-sizing: border-box; transition: box-shadow 0.28s cubic-bezier(0.4, 0, 0.2, 1) 0s; border-radius: 2px; border: none; cursor: pointer; display: inline-block; font: 500 13px / 32px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; height: 32px; margin: 0px 4px; overflow: hidden; outline: none; position: relative; text-align: center; text-transform: uppercase; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-bN97Pc { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { border-radius: 50%; left: 50%; opacity: 0; padding-bottom: 200%; position: absolute; top: 50%; transition: transform 0s linear 0.2s, opacity 0.2s ease-in 0s, -webkit-transform 0s linear 0.2s; width: 200%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ksKsZd-R5U1Nd > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { transform: translate(-50%, -50%) scale(1); opacity: 1; transition: transform 0.35s ease-out 0s, opacity 0s linear 0s, -webkit-transform 0.35s ease-out 0s; visibility: visible; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me { box-shadow: none; cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae { background-color: transparent; padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { padding: 0px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { box-shadow: rgba(0, 0, 0, 0.14) 0px 2px 2px 0px, rgba(0, 0, 0, 0.12) 0px 3px 1px -2px, rgba(0, 0, 0, 0.2) 0px 1px 5px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { box-shadow: rgba(0, 0, 0, 0.14) 0px 4px 5px 0px, rgba(0, 0, 0, 0.12) 0px 1px 10px 0px, rgba(0, 0, 0, 0.2) 0px 2px 4px -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf { background-color: rgb(66, 133, 244); color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { color: rgb(66, 133, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { color: rgba(0, 0, 0, 0.54); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915 { color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-color: rgba(66, 133, 244, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915 { background-color: rgba(255, 255, 255, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { color: rgb(51, 103, 214); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae { background-color: rgba(66, 133, 244, 0.04); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae { background-color: rgba(66, 133, 244, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae { background-color: rgba(66, 133, 244, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe { border: 1px inset rgba(0, 0, 0, 0.38); background: rgb(59, 120, 231); line-height: 30px; padding: 0px 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe { border: 1px inset rgb(66, 133, 244); line-height: 30px; padding: 0px 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe { border: 1px inset rgb(66, 133, 244); line-height: 30px; padding: 0px 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915.HB1eCd-HzV7m-LgbsSe-XpnDCe { border: 1px solid rgb(255, 255, 255); line-height: 30px; padding: 0px 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { border: none; line-height: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { padding: 0px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { background-color: rgba(0, 0, 0, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { color: rgba(0, 0, 0, 0.87); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background-color: rgba(0, 0, 0, 0.04); color: rgba(0, 0, 0, 0.54); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { color: rgba(0, 0, 0, 0.87); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background-color: rgb(255, 255, 255); color: rgba(0, 0, 0, 0.26); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915 { color: rgba(255, 255, 255, 0.3); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf { background-color: rgba(0, 0, 0, 0.12); color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(66, 133, 244, 0.32); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(66, 133, 244, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-ssJRIf > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgb(51, 103, 214); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(0, 0, 0, 0.2); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-to915 > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(255, 255, 255, 0.24); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(0, 0, 0, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); text-transform: none; border: 1px solid rgb(218, 220, 224) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-fmcmS-zTETae.HB1eCd-HzV7m-LgbsSe { color: rgb(26, 115, 232); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: normal; text-transform: none; margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(95, 99, 104); text-transform: none; border: 1px solid rgb(218, 220, 224) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-ZmdkE { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-XpnDCe { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-auswjd { border-radius: 4px; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf.HB1eCd-HzV7m-LgbsSe-OWB6Me { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(60, 64, 67); opacity: 0.38; border: 1px solid rgb(241, 243, 244) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-ZmdkE { border-radius: 4px; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { border-radius: 4px; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-XpnDCe { border-radius: 4px; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-auswjd { border-radius: 4px; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe-OWB6Me { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; border: 1px solid transparent !important; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-XpnDCe { outline: highlight solid 1px; outline-offset: -4px; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-aSvl1d-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf { color: graytext; opacity: 1; border-color: graytext; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe { display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-vhaaFf-LK5yu { border-bottom-left-radius: 0px; border-top-left-radius: 0px; margin-left: -2px; margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-vhaaFf-qwU8Me { border-bottom-right-radius: 0px; border-top-right-radius: 0px; margin-left: 0px; margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe-gk6SMd { background: rgb(225, 236, 254); z-index: 1; border: 1px solid rgb(187, 212, 251) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb [class*="docs-hc"] .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe-gk6SMd { filter: invert(100%); border-width: 0px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-gk6SMd .HB1eCd-HzV7m-LgbsSe-bN97Pc { color: rgb(25, 103, 210); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-gk6SMd.HB1eCd-HzV7m-LgbsSe-XpnDCe { background: rgb(210, 227, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-gk6SMd.HB1eCd-HzV7m-LgbsSe-XpnDCe .HB1eCd-HzV7m-LgbsSe-bN97Pc { color: rgb(24, 90, 188); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe:not([class*="docs-material-button-selected"]) { color: rgb(60, 64, 67); border-color: rgb(218, 220, 224) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe:not([class*="docs-material-button-selected"]).HB1eCd-HzV7m-LgbsSe-ZmdkE { background: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-DKlKme-LgbsSe-JNdkSc .HB1eCd-HzV7m-LgbsSe:not([class*="docs-material-button-selected"]).HB1eCd-HzV7m-LgbsSe-XpnDCe { background: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-TzA9Ye-eEGnhe { position: relative; display: inline-block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb * html .VIpgJd-TzA9Ye-eEGnhe { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :first-child + html .VIpgJd-TzA9Ye-eEGnhe { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe { background: url("//ssl.gstatic.com/editor/button-bg.png") left top repeat-x rgb(221, 221, 221); border: 0px; color: rgb(0, 0, 0); cursor: pointer; list-style: none; margin: 2px; outline: none; padding: 0px; text-decoration: none; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-style: solid; border-color: rgb(170, 170, 170); vertical-align: top; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { margin: 0px; border-width: 1px 0px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { margin: 0px -1px; border-width: 0px 1px; padding: 3px 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb * html .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { left: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb * html .VIpgJd-xl07Ob-LgbsSe-SIsrTd .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { left: -1px; right: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb * html .VIpgJd-xl07Ob-LgbsSe-SIsrTd .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { right: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :first-child + html .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { left: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :first-child + html .VIpgJd-xl07Ob-LgbsSe-SIsrTd .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { left: 1px; right: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-OWB6Me { opacity: 0.3; background-image: none !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-OWB6Me .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-OWB6Me .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-OWB6Me .VIpgJd-xl07Ob-LgbsSe-cHYyed, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-OWB6Me .VIpgJd-xl07Ob-LgbsSe-j4gsHd { color: rgb(51, 51, 51) !important; border-color: rgb(153, 153, 153) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb * html .VIpgJd-xl07Ob-LgbsSe-OWB6Me { margin: 2px 1px !important; padding: 0px 1px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :first-child + html .VIpgJd-xl07Ob-LgbsSe-OWB6Me { margin: 2px 1px !important; padding: 0px 1px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-ZmdkE .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-ZmdkE .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-color: rgb(153, 204, 255) rgb(102, 153, 238) rgb(102, 153, 238) rgb(119, 170, 255) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-FNFY6c { background-color: rgb(187, 187, 187); background-position: left bottom; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-XpnDCe .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-XpnDCe .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-color: orange; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-cHYyed { padding: 0px 4px 0px 0px; vertical-align: top; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-j4gsHd { height: 15px; width: 7px; background: url("//ssl.gstatic.com/editor/editortoolbar.png") -388px 0px no-repeat; vertical-align: top; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-qwU8Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-qwU8Me .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-qwU8Me .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-LK5yu .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-LK5yu .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { margin-left: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-LK5yu .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-left: 1px solid rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-LgbsSe-vhaaFf-LK5yu.VIpgJd-xl07Ob-LgbsSe-barxie .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-left: 1px solid rgb(221, 221, 221); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe { border-radius: 2px; cursor: default; font-size: 11px; text-align: center; white-space: nowrap; margin-right: 16px; height: 27px; line-height: 27px; min-width: 54px; outline: 0px; padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-gk6SMd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe .tk3N6e-LgbsSe-RJLb9c { margin-top: -3px; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-V67aGc { margin-left: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-roVxwc { min-width: 34px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-LK5yu.tk3N6e-LgbsSe-OWB6Me { z-index: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-barxie.tk3N6e-LgbsSe-vhaaFf-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-barxie.tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 2; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-LK5yu:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-qwU8Me:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-vhaaFf-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-vhaaFf-qwU8Me { z-index: 3; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-LK5yu { margin-left: -1px; border-bottom-left-radius: 0px; border-top-left-radius: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-vhaaFf-qwU8Me { margin-right: 0px; border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-OWB6Me:active { box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc { box-shadow: none; background-color: rgb(77, 144, 254); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(71, 135, 237))); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(53, 122, 232); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(53, 122, 232))); border: 1px solid rgb(47, 91, 183); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-JbbQac-i5vt6e { box-shadow: none; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc:active { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; background: rgb(53, 122, 232); border: 1px solid rgb(47, 91, 183); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(77, 144, 254); opacity: 0.5; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc { border-radius: 0px; border: 1px solid transparent; font-size: 13px; height: 21px; line-height: 21px; margin-right: 1px; min-width: 0px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-gk6SMd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc:active { box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc .tk3N6e-LgbsSe-RJLb9c { height: 21px; opacity: 0.55; width: 21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc .tk3N6e-LgbsSe-V67aGc { display: inline-block; margin: 0px; padding: 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-gk6SMd .tk3N6e-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-ZmdkE .tk3N6e-LgbsSe-RJLb9c { opacity: 0.9; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-OWB6Me .tk3N6e-LgbsSe-RJLb9c { opacity: 0.333; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc:focus { border: 1px solid rgb(77, 144, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e { box-shadow: none; background-color: rgb(245, 245, 245); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(245, 245, 245)), to(rgb(241, 241, 241))); color: rgb(68, 68, 68); border: 1px solid rgba(0, 0, 0, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e:active, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE:active { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background: rgb(248, 248, 248); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-gk6SMd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-gk6SMd { background-color: rgb(238, 238, 238); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e.tk3N6e-LgbsSe-barxie { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(238, 238, 238)), to(rgb(224, 224, 224))); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e:focus { border: 1px solid rgb(77, 144, 254); outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-JbbQac-i5vt6e { border: 1px solid rgba(0, 0, 0, 0.1); outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e .tk3N6e-LgbsSe-RJLb9c { opacity: 0.55; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-barxie .tk3N6e-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-gk6SMd .tk3N6e-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE .tk3N6e-LgbsSe-RJLb9c { opacity: 0.9; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me .tk3N6e-LgbsSe-RJLb9c { opacity: 0.333; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c { border-radius: 1px; background-color: rgba(255, 255, 255, 0.05); border: 1px solid rgba(155, 155, 155, 0.57); font-size: 1px; height: 11px; margin: 0px 4px 0px 1px; outline: 0px; vertical-align: text-bottom; width: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-uE9yNd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-barxie { background-color: rgba(255, 255, 255, 0.65); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px inset; border: 1px solid rgb(178, 178, 178); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-auswjd { background-color: rgb(235, 235, 235); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-XpnDCe { border: 1px solid rgb(77, 144, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-kyhDef.tk3N6e-MPu53c-XpnDCe { border: 1px solid rgba(155, 155, 155, 0.57); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-kyhDef.tk3N6e-MPu53c-OWB6Me { background-color: rgb(255, 255, 255); border: 1px solid rgb(241, 241, 241); cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-qE2ISc { height: 15px; outline: 0px; width: 15px; left: 0px; position: relative; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-uE9yNd .tk3N6e-MPu53c-qE2ISc { background: image-set(url("//ssl.gstatic.com/ui/v1/menu/checkmark-partial.png") 1x, url("//ssl.gstatic.com/ui/v1/menu/checkmark-partial_2x.png") 2x) -5px -3px no-repeat; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c-barxie .tk3N6e-MPu53c-qE2ISc { background: image-set(url("//ssl.gstatic.com/ui/v1/menu/checkmark.png") 1x, url("//ssl.gstatic.com/ui/v1/menu/checkmark_2x.png") 2x) -5px -3px no-repeat; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-TUo6Hb, .XKSfm-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { box-shadow: rgba(0, 0, 0, 0.2) 0px 4px 16px; background: padding-box rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.333); outline: 0px; position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-TUo6Hb-xJ5Hnf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-xJ5Hnf { background: rgb(255, 255, 255); left: 0px; position: absolute; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.VIpgJd-TUo6Hb-xJ5Hnf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.XKSfm-Sx9Kwc-xJ5Hnf { opacity: 0.75; }

.XKSfm-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { color: rgb(0, 0, 0); padding: 30px 42px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke { background-color: rgb(255, 255, 255); color: rgb(0, 0, 0); cursor: default; font-weight: normal; line-height: 24px; margin: 0px 0px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc { height: 11px; opacity: 0.7; padding: 17px; position: absolute; right: 0px; top: 0px; width: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc::after { content: ""; background: url("//ssl.gstatic.com/ui/v1/dialog/close-x.png"); position: absolute; height: 11px; width: 11px; right: 17px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-bN97Pc { background-color: rgb(255, 255, 255); line-height: 1.4em; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { margin-top: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button { border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(245, 245, 245)), to(rgb(241, 241, 241))); border: 1px solid rgba(0, 0, 0, 0.1); color: rgb(68, 68, 68); cursor: default; font-family: inherit; font-size: 11px; height: 29px; line-height: 27px; margin: 0px 16px 0px 0px; min-width: 72px; outline: 0px; padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button:active { background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); border: 1px solid rgb(198, 198, 198); color: rgb(51, 51, 51); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button:focus { border: 1px solid rgb(77, 144, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button[disabled] { box-shadow: none; background: none rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.05); color: rgb(184, 184, 184); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc { background-color: rgb(77, 144, 254); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(71, 135, 237))); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover { background-color: rgb(53, 122, 232); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(53, 122, 232))); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active { background-color: rgb(53, 122, 232); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(53, 122, 232))); border: 1px solid rgb(47, 91, 183); color: rgb(255, 255, 255); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus { box-shadow: rgb(255, 255, 255) 0px 0px 0px 1px inset; border: 1px solid rgba(0, 0, 0, 0); outline: rgba(0, 0, 0, 0) 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled] { box-shadow: none; background: rgb(77, 144, 254); color: rgb(255, 255, 255); opacity: 0.5; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-O0r3Gd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-McfNlf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-ostUZ { width: 512px; }

.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { border-radius: 0px; box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; transition: opacity 0.218s ease 0s; background: rgb(255, 255, 255); border: 1px solid rgba(0, 0, 0, 0.2); cursor: default; font-size: 13px; margin: 0px; outline: none; padding: 6px 0px; position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border-radius: 2px; background-color: rgb(245, 245, 245); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(245, 245, 245)), to(rgb(241, 241, 241))); border: 1px solid rgb(220, 220, 220); color: rgb(68, 68, 68); cursor: default; font-size: 11px; line-height: 27px; list-style: none; margin: 0px 2px; min-width: 46px; outline: none; padding: 0px 18px 0px 6px; text-align: center; text-decoration: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { background-color: rgb(255, 255, 255); border-color: rgb(243, 243, 243); color: rgb(184, 184, 184); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; border-color: rgb(198, 198, 198); color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { border-color: rgb(77, 144, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(238, 238, 238)), to(rgb(224, 224, 224))); border: 1px solid rgb(204, 204, 204); color: rgb(51, 51, 51); z-index: 2; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { vertical-align: top; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(119, 119, 119) transparent; border-style: solid; border-width: 4px 4px 0px; height: 0px; width: 0px; position: absolute; right: 5px; top: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c { margin-top: -3px; opacity: 0.55; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-gk6SMd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-RJLb9c { opacity: 0.9; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-gk6SMd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { border-color: rgb(89, 89, 89) transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-qwU8Me { z-index: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { z-index: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-qwU8Me:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-qwU8Me { z-index: 2; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-LK5yu:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-LK5yu { z-index: 2; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-LK5yu { margin-left: -1px; border-bottom-left-radius: 0px; border-top-left-radius: 0px; min-width: 0px; padding-left: 0px; vertical-align: top; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-vhaaFf-qwU8Me { margin-right: 0px; border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-pWKtN, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-SFgmFf { position: relative; color: rgb(51, 51, 51); cursor: pointer; list-style: none; margin: 0px; padding: 6px 8em 6px 30px; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-RDtZlf .VIpgJd-j7LFlb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-GP8zAc .VIpgJd-j7LFlb { padding-left: 16px; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-KEZkZ .VIpgJd-j7LFlb { padding-right: 44px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-x29Bmf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-bN97Pc { color: rgb(204, 204, 204) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-Bz112c { opacity: 0.3; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-ZmdkE { background-color: rgb(238, 238, 238); border-color: rgb(238, 238, 238); border-style: dotted; border-width: 1px 0px; padding-top: 5px; padding-bottom: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-ZmdkE .VIpgJd-j7LFlb-bN97Pc { color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-MPu53c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-Bz112c { background-repeat: no-repeat; height: 21px; left: 3px; position: absolute; right: auto; top: 3px; vertical-align: middle; width: 21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-wQNmvb-gk6SMd { background-image: url("//ssl.gstatic.com/ui/v1/menu/checkmark.png"); background-repeat: no-repeat; background-position: left center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-bN97Pc { color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-x29Bmf { color: rgb(119, 119, 119); direction: ltr; left: auto; padding: 0px 6px; position: absolute; right: 0px; text-align: right; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-PQTlnb-brjg8b { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-PQTlnb-hgDUwe { color: rgb(119, 119, 119); font-size: 12px; padding-left: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe { border-radius: 2px; user-select: none; background: 0px center; border-color: transparent; border-style: solid; border-width: 1px; outline: none; padding: 0px; height: 24px; color: rgb(68, 68, 68); line-height: 24px; list-style: none; text-decoration: none; vertical-align: middle; cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border: 0px; vertical-align: top; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { margin: 0px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { padding: 0px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-ZmdkE { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-gk6SMd { color: rgb(34, 34, 34); padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE { color: rgb(34, 34, 34); border-color: rgb(198, 198, 198) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { color: rgb(34, 34, 34); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-ZmdkE { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 1px; background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-auswjd { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(246, 246, 246); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(246, 246, 246)), to(rgb(241, 241, 241))); border-color: rgb(198, 198, 198); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-gk6SMd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-barxie, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-FNFY6c { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 2px inset; background-color: rgb(238, 238, 238); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(238, 238, 238)), to(rgb(224, 224, 224))); border-color: rgb(204, 204, 204); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-OWB6Me { opacity: 0.3; color: rgb(34, 34, 34) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-qwU8Me .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu .VIpgJd-INgbqf-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe-vhaaFf-LK5yu .VIpgJd-INgbqf-LgbsSe-SmKAyb-Q4BLdf { margin-left: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/ui/v1/disclosure/small-grey-disclosure-arrow-down.png") center center no-repeat; float: right; margin: 10px 2px 0px 3px; padding: 0px; opacity: 0.8; vertical-align: middle; width: 5px; height: 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-hgDUwe { border-left: 1px solid rgb(204, 204, 204); height: 17px; line-height: normal; list-style: none; margin: 0px 2px; outline: none; overflow: hidden; padding: 0px; text-decoration: none; vertical-align: middle; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-O1htCb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/ui/v1/disclosure/small-grey-disclosure-arrow-down.png") center center no-repeat; height: 11px; margin-top: 7px; width: 7px; transform: none; filter: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe-cHYyed { padding: 0px; margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar { height: 16px; overflow: visible; width: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-button { height: 0px; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track { background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 0px 0px 0px 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal { border-width: 4px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.1) 1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track:active { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.2) 1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(255, 255, 255, 0.2) 0px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-track:active { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.25) 1px 0px 0px inset, rgba(255, 255, 255, 0.15) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(255, 255, 255, 0.25) 0px 1px 0px inset, rgba(255, 255, 255, 0.15) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-thumb { background-color: rgba(0, 0, 0, 0.2); background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 1px 1px 1px 6px; min-height: 28px; padding: 100px 0px 0px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-thumb:horizontal { border-width: 6px 1px 1px; padding: 0px 0px 0px 100px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-thumb:hover { background-color: rgba(0, 0, 0, 0.4); box-shadow: rgba(0, 0, 0, 0.25) 1px 1px 1px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-thumb:active { background-color: rgba(0, 0, 0, 0.5); box-shadow: rgba(0, 0, 0, 0.35) 1px 1px 3px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-thumb { background-color: rgba(255, 255, 255, 0.3); box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-thumb:horizontal { box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-thumb:hover { background-color: rgba(255, 255, 255, 0.6); box-shadow: rgba(255, 255, 255, 0.37) 1px 1px 1px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-thumb:active { background-color: rgba(255, 255, 255, 0.75); box-shadow: rgba(255, 255, 255, 0.5) 1px 1px 3px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc::-webkit-scrollbar-track { border-width: 0px 1px 0px 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc::-webkit-scrollbar-track:horizontal { border-width: 6px 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.035); box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc-to915.tk3N6e-qrhCuc::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.07); box-shadow: rgba(255, 255, 255, 0.25) 1px 1px 0px inset, rgba(255, 255, 255, 0.15) -1px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc::-webkit-scrollbar-thumb { border-width: 0px 1px 0px 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc::-webkit-scrollbar-thumb:horizontal { border-width: 6px 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc::-webkit-scrollbar-corner { background: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body.tk3N6e-qrhCuc::-webkit-scrollbar-track-piece { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 0px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body.tk3N6e-qrhCuc::-webkit-scrollbar-track-piece:horizontal { border-width: 3px 0px 0px; box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body.tk3N6e-qrhCuc::-webkit-scrollbar-thumb { border-width: 1px 1px 1px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body.tk3N6e-qrhCuc::-webkit-scrollbar-thumb:horizontal { border-width: 5px 1px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body.tk3N6e-qrhCuc::-webkit-scrollbar-corner { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 3px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd { box-shadow: rgba(0, 0, 0, 0.2) 0px 1px 3px; background-color: rgb(255, 255, 255); border-width: 1px; border-style: solid; border-image: initial; border-color: rgb(187, 187, 187) rgb(187, 187, 187) rgb(168, 168, 168); padding: 16px; position: absolute; z-index: 1201 !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-kmh2Gb { background: url("//ssl.gstatic.com/ui/v1/icons/common/x_8px.png") no-repeat; border: 1px solid transparent; height: 21px; opacity: 0.4; outline: 0px; position: absolute; right: 2px; top: 2px; width: 21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-kmh2Gb:focus { border: 1px solid rgb(77, 144, 254); opacity: 0.8; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-hFsbo { position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { display: block; height: 0px; position: absolute; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc { border: 9px solid; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border: 8px solid; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb { bottom: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf { top: -9px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-y6n2Me { left: -9px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-cX0Lwc { right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { left: -9px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc { border-bottom-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG { border-color: rgb(255, 255, 255) transparent; left: -8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG { border-bottom-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { border-top-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG { border-top-width: 0px; top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc { border-color: transparent rgb(187, 187, 187); top: -9px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG { border-color: transparent rgb(255, 255, 255); top: -8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc { border-left-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG { border-left-width: 0px; left: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG { border-right-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc { border-radius: 0px; box-shadow: none; background-color: rgb(42, 42, 42); border: 1px solid rgb(255, 255, 255); color: rgb(255, 255, 255); cursor: default; display: block; margin-left: -1px; opacity: 1; padding: 7px 9px; position: absolute; visibility: visible; white-space: pre-wrap; word-break: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-ZYIfFd { opacity: 0; visibility: hidden; left: 20px !important; top: 20px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-wZVHld { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-hFsbo { pointer-events: none; position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { content: ""; display: block; height: 0px; position: absolute; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc { border: 6px solid; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { border: 5px solid; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-Ya1KTb { bottom: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-d6mlqf { top: -6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-y6n2Me { left: -6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-cX0Lwc { right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc { border-color: rgb(255, 255, 255) transparent; left: -6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-color: rgb(42, 42, 42) transparent; left: -5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG { border-bottom-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc { border-top-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-top-width: 0px; top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc { border-color: transparent rgb(255, 255, 255); top: -6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG { border-color: transparent rgb(42, 42, 42); top: -5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc { border-left-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG { border-left-width: 0px; left: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG { border-right-width: 0px; }

.XKSfm-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { z-index: 1001; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-xJ5Hnf { z-index: 1000; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc { background-image: none; }

.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { z-index: 2001; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb { width: 11px; height: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd { width: 11px; height: 11px; margin: auto; vertical-align: top; cursor: pointer; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd { background-color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { width: 11px; height: 11px; margin: 0px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { width: 11px; min-width: 11px; height: 11px; min-height: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb > .VIpgJd-j7LFlb { padding-left: 10px; padding-right: 10px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-KjQ5hb > .VIpgJd-j7LFlb { padding-left: 15px; padding-right: 15px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { background-color: rgb(11, 87, 208); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-barxie, .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-MPu53c.HB1eCd-HzV7m-UMrnmb-MPu53c-XpnDCe { border-color: rgb(11, 87, 208); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { color: black; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; white-space: normal; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { font-size: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe { margin: 0px 8px 0px 0px; min-width: 24px; vertical-align: middle; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-ZmdkE { box-shadow: none; background-color: rgba(0, 0, 0, 0.06); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-auswjd { box-shadow: none; background-color: rgba(0, 0, 0, 0.12); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: white; color: rgb(26, 115, 232); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(218, 220, 224) !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(241, 243, 244) !important; }

@media (forced-colors: active) {
  .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-XpnDCe { outline: highlight solid 1px; outline-offset: -4px; }
}

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(193, 216, 251) !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(204, 224, 252) !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { background: rgb(225, 236, 254); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(187, 212, 251) !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; height: 24px; padding: 3px 12px 5px; border: 1px solid transparent !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid transparent !important; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; height: 24px; padding: 3px 12px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke { font-size: 16px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb .XKSfm-Sx9Kwc-r4nke { font-size: 22px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: normal; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .lI7fHe-XKSfm.XKSfm-Sx9Kwc { width: 300px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .lI7fHe-XKSfm .XKSfm-Sx9Kwc-r4nke-fmcmS { display: block; width: 220px; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(11, 87, 208); color: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e { background: white; color: rgb(11, 87, 208); border-color: rgb(199, 199, 199) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { height: 36px; line-height: 16px; padding: 9px 16px; color: rgb(31, 31, 31); cursor: default; background: rgba(31, 31, 31, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { height: 36px; line-height: 16px; padding: 9px 16px; background-color: rgba(11, 87, 208, 0.08); box-shadow: none; color: rgb(11, 87, 208); border-color: rgb(199, 199, 199) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-auswjd { border-width: 1px; border-style: solid; border-image: initial; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background-color: rgba(11, 87, 208, 0.12); box-shadow: none; color: rgb(11, 87, 208); border-color: rgb(11, 87, 208) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(228, 228, 228); color: rgb(31, 31, 31); cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd { border: 1px solid transparent; border-radius: 100px; box-sizing: border-box; cursor: pointer; font-family: "Google Sans", Roboto, sans-serif; font-size: 14px; font-weight: 500; white-space: nowrap; height: 36px; line-height: 16px; padding: 9px 16px; background: rgb(41, 107, 214); color: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { height: 36px; line-height: 16px; padding: 9px 16px; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 2px 6px 2px; background: rgb(30, 100, 212); color: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe { background: none; border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-auswjd { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC { background-color: rgb(245, 245, 245); cursor: pointer; direction: ltr; position: relative; width: 240px; border: none; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px; border-radius: 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC { background-color: rgb(255, 255, 255); border: 1px solid rgba(60, 64, 67, 0.15); box-shadow: none; width: 282px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC { min-width: 282px; width: calc(100% - 50px); max-width: calc(50ch + 24px); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:hover { border-color: transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover { border-color: transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-k4Qmrd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC { border-radius: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC { cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:hover { background-color: transparent; cursor: pointer; border: none; box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-Nk0Zid, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-Nk0Zid .HB1eCd-Bz112c { min-height: 24px; min-width: 24px; max-width: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Nk0Zid-nUpftc.wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Nk0Zid-nUpftc.wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-Nk0Zid-nUpftc:not(.wvGCSb-pnL5fc-auswjd):hover .wvGCSb-efwuC-Nk0Zid.HB1eCd-HzV7m .HB1eCd-Bz112c .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_dark.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:active { outline: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-k4Qmrd { max-height: inherit; overflow: hidden auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-bN97Pc { overflow: hidden auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { border: none; display: none; padding: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc.wvGCSb-UbLY0d-YPqjbf-BeDmAc { padding-top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-UbLY0d-YPqjbf-BeDmAc { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd .wvGCSb-efwuC-k4Qmrd { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { display: block; height: 26px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-c6xFrd { text-align: left; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-UbLY0d-YPqjbf-BeDmAc { padding-top: 0px; border-top: none !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(119, 119, 119); font-size: 12px; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin-top: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; letter-spacing: 0.3px; line-height: 16px; }

.wvGCSb-neVct-uNfmef.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC { position: absolute; user-select: text; z-index: 500; }

.wvGCSb-neVct-uNfmef.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-CTWaPd-ZiwkRe.wvGCSb-efwuC { z-index: 502; }

.wvGCSb-neVct-uNfmef.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC { z-index: 501; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC { box-shadow: rgba(0, 0, 0, 0.2) 0px 2px 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-aIWppb { margin-right: 10px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-BvBYQ .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb.wvGCSb-JYA2rd-dHwMxe { background-color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-Bz112c-qE2ISc { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Bz112c-qE2ISc { margin-top: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-neVct-uNfmef-DF0uNb .wvGCSb-efwuC:hover { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-VkLyEc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-DyVDA { color: rgb(17, 85, 204); font-size: 11px; margin: 0px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-VkLyEc:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-DyVDA:hover { text-decoration: underline; cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-IbE0S { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-aIWppb { margin: 8px 7px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-H9tDt-xtcdFb-JIbuQc-fmcmS-sM5MNb { padding: 8px 0px 0px; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-giiMnc-GMvhG-fmcmS { overflow-wrap: break-word; margin: 8px -8px 0px; padding: 8px 8px 4px; border-color: rgb(229, 229, 229); border-top-style: solid; border-top-width: 1px; color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; line-height: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-lCdvJf-fj0AZd { background-color: rgba(140, 196, 116, 0.5); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-gk6SMd-lCdvJf-fj0AZd { background-color: rgb(140, 196, 116); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc:focus { outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe { border-top: none; border-right: none; border-left: none; border-image: initial; border-bottom: 1px solid rgb(229, 229, 229); padding: 3px 8px 5px; zoom: 1; background: rgb(245, 245, 245); position: static; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { box-shadow: rgba(0, 0, 0, 0.2) 0px 3px 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc { background-color: rgb(255, 255, 255); border-bottom: none; border-top: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe { background-color: rgb(255, 255, 255); border-bottom: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-YPqjbf-BeDmAc { background-color: rgb(255, 255, 255); border-bottom: none; border-top: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe { border-top: none; color: rgb(26, 115, 232); letter-spacing: 0.2px; margin: 0px 8px; padding: 0px; position: relative; text-align: center; -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe:not([style*="display: none"]) + .wvGCSb-Vq7Udc:not([style*="display: none"]), .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe:not([style*="display: none"]) ~ .wvGCSb-Vq7Udc[style*="display: none"] + .wvGCSb-Vq7Udc:not([style*="display: none"]) { border-top: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-Vq7Udc { padding: 8px 0px; margin: 0px 12px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { border-bottom: none; padding: 12px 12px 8px; margin: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 12px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-LgbsSe-oKdM2c { padding-top: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-bN97Pc > .wvGCSb-Vq7Udc:last-of-type, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-pnL5fc-C58Yv:only-child .wvGCSb-Vq7Udc { padding-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { padding: 8px; border-bottom: 1px solid rgb(221, 221, 221); background: rgb(255, 255, 255); min-height: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-BxnCYe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-IIEkAe .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-efwuC { background: rgb(238, 238, 238); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-yqoORe .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { border: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-YLEF4c { display: block; left: 0px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc.wvGCSb-eKrold-r08add { border-top: none !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { margin: 2px 0px 0px; color: rgb(51, 51, 51); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; font-weight: 500; height: 18px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { color: rgb(60, 64, 67); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 20px; margin-top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM .wvGCSb-Vq7Udc-FDWhSe { line-height: 1.4; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { line-height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { overflow-wrap: break-word; color: rgb(51, 51, 51); padding: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { color: rgb(0, 0, 0); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; letter-spacing: 0.2px; line-height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy { padding: 3px 21px 3px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc { background-color: rgb(241, 243, 244); border-radius: 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background: white; border-radius: 50%; bottom: -3px; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; display: flex; -webkit-box-pack: center; justify-content: center; padding: 0px; position: absolute; right: -14px; width: 32px; z-index: 10; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM a { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { margin: 0px; color: rgb(119, 119, 119); font-size: 11px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .QpLw9-qnnXGd-lI7fHe .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { -webkit-box-align: center; align-items: center; display: inline-flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb { color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; letter-spacing: 0.3px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-MGbz6c .wvGCSb-RmniWd-mQXP { -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-align: center; align-items: center; background-color: rgb(26, 115, 232); border-radius: 9px; color: white; height: 16px; -webkit-box-pack: center; justify-content: center; margin: auto 0px; overflow: hidden; transform-origin: left center; transition: transform 0.2s ease-out 0s, color 0.1s ease-in 0s, border-radius 0.2s ease 0s, -webkit-transform 0.2s ease-out 0s; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-MGbz6c:not(:hover) .wvGCSb-RmniWd-mQXP { border-radius: 50%; color: white; width: 6px; transform: scale(0.375); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc span + .wvGCSb-RmniWd-mQXP { margin-left: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-mQXP { font-weight: 600; display: inline-block; font-size: 0.75rem; font-family: Roboto, sans-serif; padding: 0px 5px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-MGbz6c:not(:hover) .wvGCSb-RmniWd-Ne3sFf { color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { min-width: 28px; width: 28px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd { height: 28px; margin: 0px; position: relative; top: auto; display: inline-block; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { height: 28px; margin: 0px; position: relative; top: auto; right: auto; display: inline-block; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd { right: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd div, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd div { margin: 1px auto auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd { border-radius: 3px 0px 0px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ERydpb-ldDtVd { border-radius: 0px 3px 3px 0px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd path, .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ERydpb-ldDtVd path { fill: rgb(26, 115, 232); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me path, .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me path { fill: rgb(60, 64, 67); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me, .wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me { background-color: white; opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd.tk3N6e-LgbsSe-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ERydpb-ldDtVd.tk3N6e-LgbsSe-OWB6Me { background-color: rgb(249, 249, 249); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC .wvGCSb-eKrold-bMcfAe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-BxnCYe .wvGCSb-eKrold-bMcfAe { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe-qAWA2 { overflow-wrap: break-word; color: rgb(17, 85, 204); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-BxnCYe-qAWA2:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2 { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:hover { text-decoration: underline; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2 { position: relative; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-BxnCYe-RWgCYc { border-top: 1px solid rgb(218, 220, 224); height: 50%; position: absolute; top: 50%; width: 100%; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd { background-color: rgb(255, 255, 255); display: inline-block; margin: 0px 20px; padding: 0px 8px; position: relative; overflow-wrap: break-word; word-break: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-rM9Gsd-eKrold { position: relative; margin: 6px 0px; padding: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-rM9Gsd-eKrold { margin-bottom: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-rM9Gsd-eKrold.wvGCSb-rM9Gsd-eKrold-xFQqWe { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold { height: 78px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 81px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-OCFbXc { color: rgb(17, 85, 204); display: none; opacity: 1; width: 100%; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-z5C9Gb:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-OCFbXc:focus { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-z5C9Gb { bottom: 0px; padding-top: 16px; position: absolute; right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { cursor: pointer; font-size: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc { background: rgb(245, 245, 245); padding: 2px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { padding: 7px 0px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-OCFbXc { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-z5C9Gb:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ti6hGc-OCFbXc:hover { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(245, 245, 245); filter: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-qAWA2-eKrold > .wvGCSb-eKrold-TJEFFc > .wvGCSb-ti6hGc-z5C9Gb { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-qAWA2-eKrold > .wvGCSb-eKrold-TJEFFc { height: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc > .wvGCSb-ti6hGc-z5C9Gb { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 100%; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc { background: rgb(245, 245, 245); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-OCFbXc { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj { margin: 6px 0px; height: 38px; white-space: nowrap; display: flex; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj { margin-top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-tJHJj { margin: 0px 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-yqoORe .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-tJHJj { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-UwkkNe { white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:hover .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-CTWaPd-ZiwkRe .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd { border: 1px solid rgba(255, 255, 255, 0.7); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .VIpgJd-xl07Ob { z-index: 600; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-UwkkNe:hover .wvGCSb-ERydpb-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-UwkkNe:hover .wvGCSb-eKrold-WlKKfd-LgbsSe { border-top-right-radius: 0px; border-bottom-right-radius: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-UwkkNe > .wvGCSb-ERydpb-ldDtVd:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-UwkkNe > .wvGCSb-eKrold-WlKKfd-LgbsSe:hover { border-top-right-radius: 2px; border-bottom-right-radius: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-UwkkNe { padding: 4px 0px 4px 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-no16zc-ldDtVd { margin-right: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-fXZhbb { padding-left: 10px; overflow: hidden; white-space: nowrap; text-overflow: ellipsis; -webkit-box-flex: 1; flex-grow: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .QpLw9-qnnXGd-lI7fHe .wvGCSb-Vq7Udc-fXZhbb span { overflow: hidden; text-overflow: ellipsis; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-fXZhbb { display: flex; -webkit-box-align: start; align-items: start; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-fXZhbb > * { overflow: hidden; text-overflow: ellipsis; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-fXZhbb > * { align-self: stretch; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { max-width: 32px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { height: 38px; margin-top: 2px; max-width: 36px; width: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { position: relative; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { margin-left: 2px; margin-top: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd { display: inline-block; margin: 0px; opacity: 0.2; position: relative; padding: 0px 4px; min-width: 50px; height: 28px; vertical-align: top; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; letter-spacing: 0.25px; line-height: 16px; background: white; color: rgb(26, 115, 232); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-WlKKfd-LgbsSe-nVMfcd:hover { background: rgb(248, 251, 255); height: 24px; padding: 3px 12px 5px; border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-WlKKfd-LgbsSe { border-radius: 3px 0px 0px 3px; display: inline-block; margin: 1px auto auto; padding: 0px; position: relative; top: auto; right: auto; vertical-align: middle; width: 28px; height: 28px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC:hover .wvGCSb-eKrold-WlKKfd-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-WlKKfd-LgbsSe { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-eKrold-DyVDA { margin-left: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-FDWhSe { overflow-wrap: break-word; color: rgb(119, 119, 119); margin: 8px -8px 0px; padding: 8px 8px 4px; border-color: rgb(229, 229, 229); border-top-style: solid; border-top-width: 1px; font-size: 11px; font-style: italic; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc-FDWhSe { color: rgb(128, 134, 139); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS { color: rgb(112, 112, 112); font-style: italic; overflow-wrap: break-word; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS { color: rgb(128, 134, 139); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; letter-spacing: 0.2px; line-height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JIbuQc-fmcmS-cGMI2b-sM5MNb { padding: 8px 0px 3px; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-Vq7Udc:last-of-type .wvGCSb-JIbuQc-fmcmS-cGMI2b-sM5MNb { padding: 8px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-GyPgRd-sM5MNb { display: flex; flex-wrap: wrap; padding-top: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border: 1px solid rgba(60, 64, 67, 0.15); border-radius: 15px; margin: 1.5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-image: radial-gradient(ghostwhite, lavender); cursor: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-eKrold-r08add.wvGCSb-Vq7Udc { padding: 16px 16px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-pnL5fc-C58Yv :only-child.wvGCSb-Vq7Udc { padding-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC { background: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(243, 246, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { border: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-k4Qmrd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd { border-radius: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-YPqjbf-BeDmAc.wvGCSb-YPqjbf .wvGCSb-YPqjbf-B7I4Od:focus { background: rgb(255, 255, 255); border: 1px solid rgb(199, 199, 199); border-radius: 18px; color: rgb(31, 31, 31); font-family: "Google Sans", Roboto, sans-serif; padding: 8px 7px 8px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { border-color: rgb(199, 199, 199); margin: 0px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-efwuC-YPqjbf-BeDmAc { border-color: rgb(199, 199, 199); margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC .wvGCSb-Vq7Udc { padding-left: 16px; padding-right: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM a { color: rgb(11, 87, 208); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(231, 237, 248); box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd.wvGCSb-efwuC:hover { background: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd:hover .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd:hover .wvGCSb-efwuC-YPqjbf-BeDmAc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-Vq7Udc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-efwuC-YPqjbf-BeDmAc { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd:hover { box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-UwkkNe { opacity: 0; transition: opacity 0.25s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-WlKKfd-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd { border: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-no16zc-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ERydpb-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-Vq7Udc-UwkkNe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-Vq7Udc-UwkkNe { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-oQLbGe { color: rgb(31, 31, 31); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-Vq7Udc-biJjHb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-biJjHb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-JIbuQc-fmcmS, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-JIbuQc-fmcmS { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; font-size: 12px; font-style: normal; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-H9tDt-xtcdFb-JIbuQc-fmcmS-sM5MNb { padding-bottom: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-no16zc-ldDtVd div, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-ERydpb-ldDtVd div { margin-top: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 0px 0px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RDNXzf-P7Vtfd .wvGCSb-efwuC-YPqjbf-BeDmAc { padding: 0px 16px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe { margin: 0px 16px; background: none; color: rgb(68, 71, 70); font: 500 14px / 20px "Google Sans", Roboto, sans-serif; -webkit-font-smoothing: antialiased; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe-qAWA2 { background: none; color: rgb(68, 71, 70); font: 500 14px / 20px "Google Sans", Roboto, sans-serif; -webkit-font-smoothing: antialiased; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd { border-radius: 100px; margin: 0px 8px; padding: 2px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(237, 242, 250); display: inline-block; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(243, 246, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd { color: rgb(11, 87, 208); text-decoration: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(231, 237, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-BxnCYe-qAWA2-k4Qmrd-haAclf { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:hover { background-color: rgba(11, 87, 208, 0.08); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-BxnCYe-qAWA2-k4Qmrd:active { background-color: rgba(11, 87, 208, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc { background-color: rgba(68, 71, 70, 0.08); border-radius: 8px; outline: transparent solid 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { box-shadow: rgba(0, 0, 0, 0.3) 0px 2px 3px, rgba(0, 0, 0, 0.15) 0px 6px 10px 4px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border-color: rgb(199, 199, 199); margin: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-XpnDCe { border-color: transparent; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 2px 6px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-color: rgb(225, 227, 225); background-image: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(237, 242, 250); font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC .wvGCSb-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb { background: rgb(243, 246, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(231, 237, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC:hover .wvGCSb-eKrold-r08add .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-efwuC.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(237, 242, 250); }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-z5C9Gb, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-ti6hGc-OCFbXc, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-pnL5fc-KUPHr-zJtgdf:hover .wvGCSb-ti6hGc-z5C9Gb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-YLEF4c-ZYyEqf { max-width: 34px; width: 34px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc-tJHJj .wvGCSb-YLEF4c { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-r08add .wvGCSb-Vq7Udc-UwkkNe { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold { height: 81px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-qAWA2-eKrold-Wz3zdc-FF2pW > .wvGCSb-eKrold-TJEFFc { height: 87px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-mQXP.wvGCSb-RmniWd-mQXP { background-color: rgb(11, 87, 208); font: 500 11px / 16px "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-ti6hGc-OCFbXc { color: rgb(11, 87, 208); text-decoration: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Vq7Udc .wvGCSb-Vq7Udc-qJTHM span, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-qJTHM .wvGCSb-eKrold-qJTHM span { color: rgb(68, 71, 70) !important; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-ZmdkE, .HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-XpnDCe { padding: 0px; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Vq7Udc .wvGCSb-lCdvJf-fj0AZd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-gk6SMd-lCdvJf-fj0AZd { background-color: highlight; color: highlighttext; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-qJTHM-Wz3zdc-ljegy-AHe6Kc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { outline: highlight solid 1px; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-itKi9e-Btuy5e-haAclf { width: fit-content; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-itKi9e-Btuy5e { cursor: pointer; display: flex; height: 18px; margin: 4px 0px 8px; outline: transparent solid 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-itKi9e-Btuy5e.HB1eCd-Guievd-WqyaDf { border: 1px solid transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-itKi9e-Btuy5e .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb docs-blue-tint-icon-cleanup .wvGCSb-itKi9e-Btuy5e .HB1eCd-HzV7m .HB1eCd-Bz112c-MqcBrc-s4vhY { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-itKi9e-Btuy5e-fmcmS { color: rgb(26, 115, 232); font: 500 14px "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e { -webkit-box-align: center; align-items: center; border-radius: 12px; height: 24px; padding: 2px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:hover { background: rgba(11, 87, 208, 0.08); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-itKi9e-Btuy5e:active { background: rgba(11, 87, 208, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId { border-bottom: 1px solid rgb(221, 221, 221); padding: 7px 10px 7px 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId { border-bottom: 1px solid rgb(218, 220, 224); padding: 12px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId { padding: 10px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId .wvGCSb-GpPaId-Bz112c-haAclf { position: absolute; right: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId table { border-spacing: 0px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-jf2N7b { background-color: rgb(242, 242, 242); color: rgb(51, 51, 51); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-jf2N7b { background-color: rgb(232, 240, 254); color: rgb(60, 64, 67); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-dHwMxe { background-color: rgb(66, 133, 244); color: white; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-dHwMxe { background-color: rgb(26, 115, 232); color: rgb(255, 255, 255); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-YLEF4c-haAclf { padding: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-YLEF4c.wvGCSb-YLEF4c { position: relative; display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-qKNFTe { padding: 0px 0px 0px 10px; width: 100%; max-width: 135px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-V67aGc { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; letter-spacing: 0.3px; line-height: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-V67aGc { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-JYA2rd-fmcmS { font-weight: 500; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId-JYA2rd-fmcmS { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; letter-spacing: 0.25px; line-height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-Bz112c-qE2ISc-JaPV2b { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-Bz112c-qE2ISc-HLvlvd { margin-top: 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-Bz112c-qE2ISc-HLvlvd { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe { width: 28px; height: 28px; min-width: 28px; padding: 0px; margin: 0px; background: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe-JaPV2b { opacity: 0.2; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe-JaPV2b { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd { border: 1px solid rgba(255, 255, 255, 0.38); opacity: 0.7; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd:hover { border: 1px solid rgb(255, 255, 255); opacity: 1; background: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe-HLvlvd { border: none; opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-dhWRR-xCiRjb { margin: -15px -15px 0px; padding-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId { -webkit-box-align: center; align-items: center; border: none; box-sizing: border-box; border-radius: 4px; display: flex; -webkit-box-pack: justify; justify-content: space-between; margin: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId.wvGCSb-JYA2rd-jf2N7b { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId.wvGCSb-JYA2rd-dHwMxe .wvGCSb-GpPaId-JYA2rd-fmcmS { text-transform: uppercase; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId-V67aGc { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; line-height: 20px; letter-spacing: 0.25px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId-JYA2rd-fmcmS { margin-left: 4px; max-width: 195px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-SYOSDb-iib5kc-LgbsSe { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId { border: none; padding: 1px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId-qKNFTe { -webkit-box-align: center; align-items: center; display: flex; height: 38px; max-width: 210px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-dHwMxe { background-color: rgb(211, 227, 253); color: rgb(4, 30, 73); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-jf2N7b { background-color: inherit; color: rgb(68, 71, 70); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId-V67aGc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId-JYA2rd-fmcmS { display: inline-block; font: 500 12px / 16px "Google Sans", Roboto, sans-serif; vertical-align: middle; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId-V67aGc { font: 500 12px / 16px "Google Sans", Roboto, sans-serif; vertical-align: middle; white-space: nowrap; display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId-JYA2rd-fmcmS { margin: 0px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId .wvGCSb-Bz112c-qE2ISc-JaPV2b { margin-top: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe { background: none; border-radius: 100%; height: 32px; width: 32px; margin: 0px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-GpPaId .wvGCSb-SYOSDb-iib5kc-LgbsSe.tk3N6e-LgbsSe-auswjd { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId .wvGCSb-GpPaId-Bz112c-haAclf { right: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-dhWRR-xCiRjb { padding-bottom: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-JYA2rd-dHwMxe .wvGCSb-SYOSDb-iib5kc-LgbsSe .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .wvGCSb-JYA2rd-dHwMxe .wvGCSb-SYOSDb-iib5kc-LgbsSe .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(12%) sepia(17%) saturate(6039%) hue-rotate(199deg) brightness(93%) contrast(106%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-JYA2rd-jf2N7b .wvGCSb-SYOSDb-iib5kc-LgbsSe .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg"); left: -52px; top: -556px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC.wvGCSb-pnL5fc-auswjd .wvGCSb-JYA2rd-jf2N7b .wvGCSb-SYOSDb-iib5kc-LgbsSe .HB1eCd-Bz112c-RJLb9c { left: -52px; top: -9808px; }

.HB1eCd-MqDS2b-uoC0bf.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GpPaId.wvGCSb-JYA2rd-dHwMxe .wvGCSb-GpPaId-JYA2rd-fmcmS { text-transform: lowercase; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .wvGCSb-GpPaId td:last-child { text-align: end; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MwUX8 { -webkit-box-align: center; align-items: center; background-color: rgb(249, 249, 249); border: 0.0625em solid rgb(186, 186, 186); border-radius: 0.2em; bottom: 0.1em; box-sizing: border-box; display: inline-flex; height: 1.1em; -webkit-box-pack: center; justify-content: center; margin-left: 0.3em; position: relative; width: 1.8em; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .DQD9Vb { color: rgb(186, 186, 186); font-size: 0.6em; font-weight: bold; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .G337pd { color: rgb(128, 134, 139) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd { background: rgb(255, 255, 255); border: 1px solid rgb(200, 200, 200); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin: 0px; padding: 4px 0px; position: absolute; z-index: 900; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd { border-color: transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; padding: 9px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd div { cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd .ztA2jd-oKdM2c { height: auto; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd .ztA2jd-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd div.auswjd { background-color: rgb(238, 238, 238); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd .ztA2jd-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd div.auswjd { background-color: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd-AHUcCb { font-weight: bold; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-wTehdb-ORHb { background-color: rgb(254, 247, 224); padding: 8px 0px 8px 14px; margin: 12px 0px 8px; display: flex; -webkit-box-align: center; align-items: center; outline: transparent solid 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-wTehdb-ORHb { left: -12px; width: 268px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-wTehdb-ORHb { left: -8px; width: 226px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC .wvGCSb-wTehdb-ORHb-haAclf { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; width: calc(100% + 24px); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC .wvGCSb-wTehdb-ORHb { width: calc(100% - 12px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-F6aDIf.wvGCSb-wTehdb-ORHb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-F6aDIf.wvGCSb-wTehdb-ORHb { border-radius: 4px; left: 0px; width: inherit; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-efwuC .wvGCSb-F6aDIf.wvGCSb-wTehdb-ORHb { width: calc(100% - 36px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-wTehdb-ORHb { left: -56px; width: 281px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-F6aDIf.wvGCSb-wTehdb-ORHb { border-radius: 4px; left: 0px; width: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-Bz112c-SxQuSe { width: 18px; height: 18px; margin: 1px 2px 2px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb .tk3N6e-LgbsSe.wTehdb-ORHb-Tswv1b { margin-right: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .tk3N6e-LgbsSe.wTehdb-ORHb-Tswv1b { margin-left: auto; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-wTehdb-ORHb-fmcmS { font-size: 12px; width: 195px; padding-left: 10px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-neVct-uNfmef-XHgP6b-m3mY0d .wvGCSb-wTehdb-ORHb-fmcmS { width: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-wTehdb-ORHb-fmcmS { font-size: 12px; width: 188px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-wTehdb-ORHb-fmcmS { width: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-wTehdb-ORHb .tk3N6e-LgbsSe-n2to0e { min-width: 21px; padding: 0px 2px; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe.wTehdb-ORHb-Tswv1b { margin-right: 10px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { min-width: 464px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke, .wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-bN97Pc { padding-bottom: 0px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-h9d3hd { cursor: pointer; float: right; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-Dzid5 { color: rgb(95, 99, 104); font: 14px / 20px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; margin-bottom: 16px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-oKdM2c { padding-bottom: 12px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-xJzy8c { border-radius: 50%; float: left; height: 32px; margin-right: 16px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-V1ur5d { color: rgb(60, 64, 67); font: 14px / 20px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; letter-spacing: 0.2px; }

.wTehdb-MZArnb-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wTehdb-MZArnb-jOfkMb { color: rgb(95, 99, 104); font: 12px / 16px Roboto, RobotoDraft, Helvetica, Arial, sans-serif; letter-spacing: 0.3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YLEF4c { left: 0px; position: absolute; object-fit: cover; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YLEF4c { border-radius: 50%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YLEF4c-ExtcI { opacity: 0.4; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YLEF4c-ExtcI { background-color: white; opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eLiUMc-Tswv1b { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(187, 187, 187); text-align: right; padding-right: 30px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eLiUMc-Tswv1b a { color: rgb(187, 187, 187); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd { min-height: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-haAclf { background: rgb(242, 242, 242); padding: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-haAclf { background: white; padding: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-tJHJj-HiaYvf { max-width: 100%; margin-bottom: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-aAmChf-EfADOe .wvGCSb-AQdXhd-tJHJj-HiaYvf { border: 1px solid rgb(218, 220, 224); box-sizing: border-box; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-tJHJj { -webkit-box-align: center; align-items: center; color: rgb(60, 64, 67); display: flex; line-height: 20px; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; vertical-align: top; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-qAJZhe-RFnRab .wvGCSb-AQdXhd-tJHJj { color: rgb(32, 33, 36); font-size: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-aAmChf-EfADOe .wvGCSb-AQdXhd-tJHJj { color: rgb(32, 33, 36); line-height: 28px; font-size: 22px; font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-tJHJj-Bz112c { left: -3px; margin-right: 3px; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .HB1eCd-Bz112c.wvGCSb-AQdXhd-tJHJj-Bz112c-haAclf { height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-qJTHM { padding: 12px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-qAJZhe-RFnRab .wvGCSb-AQdXhd-qJTHM { color: rgb(60, 64, 67); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-qAJZhe-RFnRab-AR1m8c-wt8N5c .wvGCSb-AQdXhd-qJTHM a { display: inline-block; font-size: 14px; line-height: 20px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .stjqE-Fi6iz-qAJZhe-RFnRab-AR1m8c-wt8N5c .wvGCSb-AQdXhd-rM9Gsd { font-size: 0px; line-height: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-rM9Gsd { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; line-height: 20px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-qJTHM a { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-MPu53c-haAclf { border-bottom: 1px solid rgb(218, 220, 224); margin-bottom: 16px; padding-bottom: 16px; padding-top: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-MPu53c-haAclf .HB1eCd-HzV7m-UMrnmb-MPu53c { cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-kv69tf-ti6hGc-oFshpd-MPu53c { margin-bottom: 10px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-kv69tf-ti6hGc-oFshpd-V67aGc { color: rgb(60, 64, 67); padding-left: 10px; position: relative; top: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-ti6hGc-OCFbXc { color: rgb(17, 85, 204); cursor: pointer; font-size: 11px; outline: none; padding-top: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-ti6hGc-z5C9Gb:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-ti6hGc-OCFbXc:hover { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-c6xFrd-Ne3sFf-fmcmS { font-size: 12px; line-height: 16px; margin-bottom: 10px; padding-right: 10px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-fmcmS-zTETae-c6xFrd-haAclf { display: flex; -webkit-box-pack: end; justify-content: flex-end; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-AQdXhd-fmcmS-zTETae-c6xFrd-haAclf div.HB1eCd-HzV7m-LgbsSe { margin-left: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd { background: rgb(253, 252, 251); border: 1px solid rgb(196, 199, 197); border-radius: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd .wvGCSb-AQdXhd { border: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-haAclf { background: rgb(253, 252, 251); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:hover .wvGCSb-AQdXhd-haAclf { background: rgba(31, 31, 31, 0.08); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-efwuC:active .wvGCSb-AQdXhd-haAclf { background: rgba(31, 31, 31, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd .wvGCSb-AQdXhd-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd:hover .wvGCSb-AQdXhd-haAclf { background: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-qJTHM, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-ti6hGc-z5C9Gb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-ti6hGc-OCFbXc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-kv69tf-ti6hGc-oFshpd-V67aGc { color: rgb(68, 71, 70); font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-AQdXhd-qJTHM a { color: rgb(11, 87, 208); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c { height: 32px; color: rgb(0, 0, 0); padding: 4px 8px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c { height: 36px; padding: 6px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c .wvGCSb-YLEF4c { float: left; left: auto; position: relative; padding-right: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c .wvGCSb-YLEF4c { padding-right: 0px; margin-right: 8px; margin-top: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c-V1ur5d { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c-xvr5H { text-overflow: ellipsis; white-space: nowrap; overflow: hidden; color: rgb(119, 119, 119); font-size: 0.9em; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c-V1ur5d { color: rgb(60, 64, 67); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; line-height: 20px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-ztA2jd-AHUcCb { font-weight: 700; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-M7sy3e-oKdM2c-xvr5H { color: rgb(60, 64, 67); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; }

.wvGCSb-VkLyEc-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { font-size: 14px; white-space: normal; width: 472px; }

.wvGCSb-VkLyEc-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-VkLyEc-Sx9Kwc-VdSJob { width: 424px; }

.wvGCSb-VkLyEc-Sx9Kwc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-LgbsSe-bN97Pc { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yqoORe-Wz3zdc-Z7HxEc-nUpftc.wvGCSb-efwuC { border: unset; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; background: unset; border-radius: 24px; width: 282px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yqoORe-Wz3zdc-Z7HxEc-nUpftc-aIWppb { width: 282px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yqoORe-Wz3zdc-nKQ6qf-bEDTcc-OiiCO { animation-duration: 0.3s; animation-name: draft-emoji-slide-in; animation-timing-function: ease-in-out; animation-iteration-count: 1; }

@keyframes draft-emoji-slide-in { 
  0% { width: 20%; opacity: 0; }
}

@-webkit-keyframes draft-emoji-slide-in { 
  0% { width: 20%; opacity: 0; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { display: flex; -webkit-box-align: center; align-items: center; height: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { background-size: contain; height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { font-family: "Noto Color Emoji", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 20px; height: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-NnAfwf { -webkit-box-align: center; align-items: center; display: flex; font-size: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c-haAclf { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf > * { padding: 0px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-dIxMhd-Ca9lu.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { color: rgb(26, 115, 232); font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :not(.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-dIxMhd-Ca9lu).HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf { color: rgb(95, 99, 104); font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-PrY1nf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c-haAclf { font-size: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc { background-color: rgb(255, 255, 255); border-radius: 8px; box-shadow: rgb(189, 193, 198) 1px 0px 8px 1px; color: rgb(95, 99, 104); display: flex; font-size: 13px; font-weight: 400; line-height: 20px; margin-top: 7px; max-width: 258px; padding: 4px; text-align: center; width: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG { border-color: rgb(255, 255, 255) transparent; left: -6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { height: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb.HB1eCd-HzV7m-LgbsSe { height: 24px; padding: 0px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c { height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Bz112c.wvGCSb-Wz3zdc-gmhCAd-LgbsSe-Wz3zdc-sLO9V-qnnXGd { font-size: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-aIWppb .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-haAclf > * { padding: 0px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC { background: unset; border: unset; border-radius: 15px; max-width: 282px; width: fit-content; min-width: auto; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC:hover { box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-pnL5fc-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-pnL5fc-auswjd:hover { box-shadow: unset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd { border: 1px solid rgba(60, 64, 67, 0.15); border-radius: 15px; height: fit-content; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-qN5Z7b-LgbsSe .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd:not(:hover) { border-color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd :not(.HB1eCd-HzV7m-LgbsSe-XpnDCe).HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border-color: transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .VIpgJd-haAclf-DKlKme { display: flex; flex-wrap: wrap; -webkit-box-pack: center; justify-content: center; margin: 1.5px; max-width: 200px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-color: rgb(255, 255, 255); border: 1px solid rgba(60, 64, 67, 0.15); display: flex; border-radius: 15px; margin: 1.5px; opacity: 0; width: fit-content; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-image: radial-gradient(ghostwhite, lavender); cursor: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background-color: rgb(232, 240, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; line-height: 32px; padding: 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { padding: 1px 9px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-haAclf { display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-nK2kYb { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: reverse; flex-direction: row-reverse; -webkit-box-pack: justify; justify-content: space-between; padding: 0px 4px; margin-top: 4px; gap: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background-color: rgb(255, 255, 255); color: rgba(0, 0, 0, 0.26); border-radius: 16px; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; display: flex; -webkit-box-pack: center; justify-content: center; height: 32px; margin: 0px; padding: 0px; width: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-OWB6Me.HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { background-color: rgba(0, 0, 0, 0.04); color: rgba(0, 0, 0, 0.54); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .VIpgJd-haAclf-DKlKme { border: none; margin: 0px; gap: 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd { border: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .wvGCSb-efwuC-k4Qmrd { overflow: visible; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-efwuC:hover { background: none; box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-NnAfwf { font-family: "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-dIxMhd-Ca9lu .wvGCSb-Wz3zdc-gmhCAd-LgbsSe-NnAfwf { color: rgb(11, 87, 208); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { border: none; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf { background: rgb(243, 246, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd.wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-bN97Pc { background: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-bN97Pc { height: 100%; padding: 0px 8px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-nK2kYb { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-ZmdkE .HB1eCd-HzV7m-LgbsSe-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-ZmdkE .HB1eCd-HzV7m-LgbsSe-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf:hover .HB1eCd-HzV7m-LgbsSe-bN97Pc { background: rgba(11, 87, 208, 0.08); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-Wz3zdc-nK2kYb .HB1eCd-HzV7m-LgbsSe-XpnDCe .HB1eCd-HzV7m-LgbsSe-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe:active .HB1eCd-HzV7m-LgbsSe-bN97Pc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd.wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-XpnDCe .HB1eCd-HzV7m-LgbsSe-bN97Pc { background: rgba(11, 87, 208, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc-GyPgRd .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae { border: none; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc.wvGCSb-pnL5fc .HB1eCd-HzV7m-LgbsSe-Kb3HCc-ssJRIf:active, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae.HB1eCd-HzV7m-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae.HB1eCd-HzV7m-LgbsSe-XpnDCe { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-auswjd .HB1eCd-HzV7m-LgbsSe-MV7yeb-zTETae .HB1eCd-Bz112c { margin: 0px 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-eKrold-GyPgRd-sM5MNb .wvGCSb-Wz3zdc-Z7HxEc-lI7fHe-nUpftc .HB1eCd-HzV7m-LgbsSe-OWB6Me .HB1eCd-HzV7m-LgbsSe-bN97Pc { background-color: rgb(225, 227, 225); background-image: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c { overflow: hidden; vertical-align: middle; user-select: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/d-icons31.png"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RJLb9c-ws0Ijb::before { transform: scale(0.5); transform-origin: 0px 0px; display: inline-block; image-rendering: -webkit-optimize-contrast; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RJLb9c { }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RJLb9c-haAclf { position: absolute; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-PFprWc-JaPV2b { top: -88px; left: -4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-PFprWc-nllRtd { top: -106px; left: -4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-PFprWc-SxQuSe { height: 18px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-HzFBSb { top: -25px; left: -25px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-HzFBSb-SxQuSe { height: 13px; width: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-Ge5tnd-jNm5if { top: -48px; left: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-JaPV2b { left: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-HLvlvd { top: -140px; left: -49px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-SxQuSe { height: 21px; width: 21px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-JaPV2b { left: -42px; top: -24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-HLvlvd { top: 0px; left: -42px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-SxQuSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb .wvGCSb-Bz112c-no16zc-qE2ISc-SxQuSe { height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-ERydpb-ldDtVd-AZ4Tub { top: -44px; left: -21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-ERydpb-ldDtVd-AZ4Tub-SxQuSe { height: 21px; width: 21px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-ERydpb-ldDtVd-AZ4Tub-SxQuSe { height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-Ge5tnd-jNm5if-SxQuSe { height: 14px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RPzgNd-vfifzc-RxYbNe { left: -25px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RPzgNd-vfifzc-RxYbNe-SxQuSe { height: 21px; width: 14px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RPzgNd-vfifzc-RxYbNe { left: 0px; top: -164px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-Bz112c-RPzgNd-vfifzc-RxYbNe { top: -165px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-RPzgNd-vfifzc-RxYbNe-SxQuSe { height: 24px; width: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-hdBvUb { top: -64px; left: -2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-hdBvUb-SxQuSe { height: 21px; width: 21px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Guievd-WqyaDf .wvGCSb-Bz112c-RJLb9c { filter: invert(100%); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-DfC5c-wvGCSb-i3jM8c { top: -48px; left: 12px; height: 14px; width: 18px; position: absolute; clip: rect(48px, 20px, 72px, 0px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-DfC5c-wvGCSb-SIsrTd { top: -48px; left: 60px; height: 14px; width: 18px; position: absolute; clip: rect(48px, -28px, 63px, -48px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Guievd-WqyaDf .tk3N6e-MPu53c-barxie .tk3N6e-MPu53c-qE2ISc::before { content: url("//ssl.gstatic.com/docs/common/d-icons31.png"); position: absolute; left: -50px; top: -124px; width: 15px; height: 15px; clip: rect(125px, 65px, 140px, 51px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m > .wvGCSb-RmniWd-jNm5if-Bz112c > .wvGCSb-Bz112c-htvI8d-jNm5if { top: -125px; left: -4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m > .wvGCSb-Bz112c-htvI8d-jNm5if-SxQuSe { height: 18px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .wvGCSb-Bz112c-DfC5c-wvGCSb-i3jM8c { top: -125px; left: 11px; height: 18px; width: 18px; clip: rect(125px, 20px, 145px, 0px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m .wvGCSb-Bz112c-DfC5c-wvGCSb-SIsrTd { top: -125px; left: 59px; height: 18px; width: 18px; clip: rect(125px, -28px, 145px, -48px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-OWB6Me .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ldDtVd-LgbsSe.tk3N6e-LgbsSe-OWB6Me .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-TvD9Pc { top: -364px; left: -30px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-TvD9Pc-SxQuSe { height: 18px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-Tswv1b { top: -364px; left: -48px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Bz112c-Tswv1b-SxQuSe { height: 18px; width: 18px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye .HB1eCd-ldDtVd-LgbsSe:not(.tk3N6e-LgbsSe-OWB6Me) .HB1eCd-HzV7m .HB1eCd-Bz112c-RJLb9c::before { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf { position: relative; outline: none; zoom: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf.wvGCSb-YPqjbf-mOyJmb { display: block !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lvBGLe { cursor: text; text-align: start; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lvBGLe:empty::before { color: rgb(128, 134, 139); content: attr(placeholder); display: block; pointer-events: none; }

@media screen and (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lvBGLe:empty::before { color: graytext; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lvBGLe p { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-B7I4Od { box-sizing: border-box; color: rgb(153, 153, 153); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 13px; margin: 0px; overflow: hidden; padding: 4px; resize: none; width: 100%; border: 1px solid rgb(200, 200, 200); outline-width: 0px !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-B7I4Od { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(60, 64, 67); font-size: 14px; line-height: 20px; min-height: 36px; padding: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-B7I4Od:focus { border: 2px solid rgb(26, 115, 232); box-shadow: none; padding: 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-B7I4Od:disabled { background-color: rgb(238, 238, 238) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :first-child + html .wvGCSb-YPqjbf-B7I4Od { width: 95%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-c6xFrd { display: none; zoom: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-c6xFrd-aIWppb { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { color: rgb(0, 0, 0); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { color: rgb(60, 64, 67); }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-B7I4Od { background-color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-YsTx5 > .wvGCSb-YPqjbf-c6xFrd { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-IIyL0-wcotoc-fmcmS { color: rgb(97, 97, 97); font-style: italic; padding: 5px 0px 3px; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b { padding: 6px 8px 4px; background-color: rgb(245, 245, 245); border-style: solid; border-width: 0px 1px 1px; border-color: rgb(200, 200, 200); margin-bottom: 8px; cursor: pointer; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b { padding: 6px 8px 11px 0px; background-color: rgb(255, 255, 255); border-width: 1px; border-style: solid; border-color: transparent transparent rgb(218, 220, 224); border-image: initial; margin-bottom: 18px; cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-Q4BLdf { margin: 2px 10px 0px 0px; float: left; width: 11px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-JYA2rd-fmcmS { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-fmcmS { text-align: left; white-space: nowrap; overflow: hidden; text-overflow: ellipsis; font-size: 13px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(112, 112, 112); font-weight: normal; display: inline-block; width: calc(100% - 51px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-fmcmS.wvGCSb-YPqjbf-JYA2rd-fmcmS-di8rgd-Q8Kwad { width: calc(100% - 23px); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-fmcmS { margin-top: 6px; margin-left: 8px; white-space: nowrap; overflow: hidden; text-overflow: ellipsis; font-size: 14px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; color: rgb(60, 64, 67); font-weight: normal; display: inline-block; width: calc(100% - 57px); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-fmcmS.wvGCSb-YPqjbf-JYA2rd-fmcmS-di8rgd-Q8Kwad { width: calc(100% - 29px); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-YPqjbf-JYA2rd-O1htCb { margin-top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JYA2rd-O1htCb-AHmuwe { border-radius: 2px; border: 1px solid rgb(77, 144, 254) !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-O1htCb { border: none; background: none; box-shadow: none; cursor: pointer; float: right; width: 24px; height: 15px; margin: 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-YPqjbf-JYA2rd-O1htCb { margin-top: 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-O1htCb .VIpgJd-xl07Ob-LgbsSe-cHYyed { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-JYA2rd-O1htCb .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JYA2rd-O1htCb-ibnC6b { padding: 0px; border-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JYA2rd-O1htCb-ibnC6b.VIpgJd-j7LFlb-sn54Q { background-color: rgb(242, 242, 242); }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.wvGCSb-JYA2rd-O1htCb-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { padding: 4px 0px; max-height: 222px; overflow-y: auto; box-sizing: border-box; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { padding: 8px 0px; }

.VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JYA2rd-O1htCb-ibnC6b, .VIpgJd-xl07Ob.VIpgJd-xl07Ob-BvBYQ.HB1eCd-UMrnmb.wvGCSb-JYA2rd-O1htCb-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-JYA2rd-O1htCb-ibnC6b.VIpgJd-xl07Ob-ibnC6b-sn54Q { border: none; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-j4gsHd { width: 24px; background: url("//ssl.gstatic.com/images/icons/material/system/2x/arrow_drop_down_black_24dp.png") center center / 24px no-repeat; opacity: 0.54; box-sizing: border-box; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-j4gsHd:hover { opacity: 0.87; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-n0tgWb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-lQVAed-b0t70b .VIpgJd-xl07Ob-LgbsSe-SmKAyb-Q4BLdf { border-style: none; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf-lvBGLe:empty::before { color: rgb(68, 71, 70); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-YPqjbf-lQVAed-b0t70b { background-color: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-aZ2wEe { height: 100px; overflow: hidden; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vyDMJf-aZ2wEe { height: 28px; left: 50%; margin-left: -14px; position: absolute; top: 36px; width: 28px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .docos-mention { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .docos-mention-current-user { -webkit-box-align: center; align-items: center; background-color: rgb(210, 227, 252); border-radius: 4px; color: rgb(23, 78, 166); padding: 2px 4px; top: 0px; width: max-content; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-H6MApb a.docos-mention-current-user { background: rgb(26, 115, 232); color: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u { background-color: rgb(255, 255, 255); border-bottom: none; border-top: 1px solid rgb(218, 220, 224); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: auto; padding: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-c6xFrd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: justify; justify-content: space-between; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe { background-image: none; border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; -webkit-box-align: center; align-items: center; color: rgb(13, 101, 45); cursor: pointer; display: flex; margin: 0px; padding: 8px; text-transform: none; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-ZmdkE { background: rgba(24, 128, 56, 0.04); color: rgb(13, 101, 45); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe { background: rgba(24, 128, 56, 0.12); color: rgb(13, 101, 45); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-auswjd { background: rgba(24, 128, 56, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-di8rgd-AHmuwe-VtOx3e { line-height: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { background-color: rgba(52, 168, 83, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-LzZ0g { -webkit-box-align: center; align-items: center; display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-MYFTse, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-tJiF1e { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-MYFTse .HB1eCd-Bz112c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-tJiF1e .HB1eCd-Bz112c { left: -3px; margin: 0px; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-MYFTse:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-tJiF1e:hover { background: rgba(32, 33, 36, 0.04); cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-MYFTse:focus, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-tJiF1e:focus { background: rgba(32, 33, 36, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-MYFTse:active, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yXBf7b-ZMv3u-tJiF1e:active { background: rgba(32, 33, 36, 0.1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-yXBf7b-ZMv3u { background: rgb(243, 246, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-KX2r4e:hover .wvGCSb-yXBf7b-ZMv3u, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-KX2r4e-auswjd .wvGCSb-yXBf7b-ZMv3u { background: rgb(231, 237, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-KX2r4e:hover .wvGCSb-yXBf7b-ZMv3u, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-qJTHM-aAmChf .wvGCSb-KX2r4e-auswjd .wvGCSb-yXBf7b-ZMv3u { background: rgb(237, 242, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe { border-radius: 100px; color: rgb(11, 87, 208); padding: 10px 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-ZmdkE { background: rgba(11, 87, 208, 0.08); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe.HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-auswjd { background: rgba(11, 87, 208, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-FNFY6c-NkyfNe-RDNXzf-LgbsSe > .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u-LzZ0g .HB1eCd-HzV7m-LgbsSe { background: none; border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u-LzZ0g .HB1eCd-HzV7m-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u-LzZ0g .HB1eCd-HzV7m-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u-LzZ0g .HB1eCd-HzV7m-LgbsSe-auswjd { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-yXBf7b-ZMv3u-LzZ0g .HB1eCd-HzV7m-LgbsSe .HB1eCd-Bz112c { left: -5px; top: -4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-bN97Pc { width: 500px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-V67aGc { padding: 0px 3px 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-bMcfAe { padding-left: 3px; margin-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-tJHJj { font-weight: 500; margin-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-h9d3hd { position: absolute; right: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb { display: inline-block; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd { background: none; border-radius: 100%; height: 32px; width: 32px; -webkit-box-align: center; align-items: center; cursor: pointer; display: flex; -webkit-box-pack: center; justify-content: center; left: -1px; margin: auto; position: relative; transition: opacity 0.25s cubic-bezier(0.4, 0, 0.2, 1) 0s; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd:hover { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; box-shadow: none; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd:focus { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; box-shadow: none; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-SmKAyb-Q4BLdf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .wvGCSb-Bz112c { margin-top: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-j4gsHd { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb .VIpgJd-j7LFlb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb.VIpgJd-xl07Ob .VIpgJd-j7LFlb { padding-right: 15px; padding-left: 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd { animation: 1568ms linear 0s infinite normal none running container-rotate; }

@-webkit-keyframes container-rotate { 
  100% { transform: rotate(1turn); }
}

@keyframes container-rotate { 
  100% { transform: rotate(1turn); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-pbTTYe { position: absolute; width: 100%; height: 100%; opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-v3pZbf { border-color: rgb(66, 133, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-oq6NAc { border-color: rgb(219, 68, 55); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-gS7Ybc { border-color: rgb(244, 180, 0); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-nllRtd { border-color: rgb(15, 157, 88); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-v3pZbf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running blue-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-oq6NAc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running red-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-gS7Ybc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running yellow-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-nllRtd { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running green-fade-in-out; }

@-webkit-keyframes fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@keyframes fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@-webkit-keyframes blue-fade-in-out { 
  0% { opacity: 1; }
  25% { opacity: 1; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 1; }
  100% { opacity: 1; }
}

@keyframes blue-fade-in-out { 
  0% { opacity: 1; }
  25% { opacity: 1; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 1; }
  100% { opacity: 1; }
}

@-webkit-keyframes red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 1; }
  50% { opacity: 1; }
  51% { opacity: 0; }
}

@keyframes red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 1; }
  50% { opacity: 1; }
  51% { opacity: 0; }
}

@-webkit-keyframes yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 1; }
  75% { opacity: 1; }
  76% { opacity: 0; }
}

@keyframes yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 1; }
  75% { opacity: 1; }
  76% { opacity: 0; }
}

@-webkit-keyframes green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 1; }
  90% { opacity: 1; }
  100% { opacity: 0; }
}

@keyframes green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 1; }
  90% { opacity: 1; }
  100% { opacity: 0; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-pehrl-TpMipd { position: absolute; box-sizing: border-box; top: 0px; left: 45%; width: 10%; height: 100%; overflow: hidden; border-color: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-pehrl-TpMipd .aZ2wEe-LkdAo { width: 1000%; left: -450%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-LkdAo-e9ayKc { display: inline-block; position: relative; width: 50%; height: 100%; overflow: hidden; border-color: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-LkdAo-e9ayKc .aZ2wEe-LkdAo { width: 200%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-LkdAo { box-sizing: border-box; height: 100%; border-width: 3px; border-style: solid; border-top-color: inherit; border-right-color: inherit; border-left-color: inherit; border-radius: 50%; animation: 0s ease 0s 1 normal none running none; border-bottom-color: transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { transform: rotate(129deg); border-right-color: transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { left: -100%; transform: rotate(-129deg); border-left-color: transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running left-spin; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running right-spin; }

@-webkit-keyframes left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@keyframes left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@-webkit-keyframes right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@keyframes right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aZ2wEe-hj4D6d { position: absolute; inset: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vyDMJf-aZ2wEe.auswjd { animation: 1568ms linear 0s infinite normal none running container-rotate; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-pbTTYe.aZ2wEe-v3pZbf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running blue-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-pbTTYe.aZ2wEe-oq6NAc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running red-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-pbTTYe.aZ2wEe-gS7Ybc { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running yellow-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-pbTTYe.aZ2wEe-nllRtd { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running green-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running left-spin; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running right-spin; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-iQd6Fc .ZYIfFd-IT5dJd-iQd6Fc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ti6hGc-IT5dJd-iQd6Fc { display: none !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-iQd6Fc .ti6hGc-IT5dJd-iQd6Fc { display: inline-block !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-WlKKfd-sn54Q { border: 1px solid rgba(0, 0, 0, 0.2); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-WlKKfd-OiiCO { transition: all 0.27s ease-out 0s; transform: scale(0.3); transform-origin: center top; opacity: 0.3; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow-wrapper { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow { background: rgba(0, 0, 0, 0.7); color: rgb(255, 255, 255); position: absolute; z-index: 700; left: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-bnBfGc-BPrWId > :focus { outline: transparent solid 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-bnBfGc-jyrRxf { height: 100%; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow-description { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow-confirm, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docos-shadow-delete { margin: 2px 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf #docos-shadow .tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf #docos-shadow .tk3N6e-LgbsSe-XpnDCe { background: white; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F9IAbd-xtcdFb { display: flex; -webkit-box-pack: justify; justify-content: space-between; text-align: center; margin-right: 6px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F9IAbd-xtcdFb-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe { -webkit-box-align: center; align-items: center; display: flex; height: auto; -webkit-box-pack: center; justify-content: center; padding: 3px 12px; white-space: normal; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F9IAbd-xtcdFb .wvGCSb-F9IAbd-xtcdFb-LgbsSe:last-child { margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F9IAbd-xtcdFb-LgbsSe-cHYyed { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb.HB1eCd-UMrnmb .wvGCSb-F9IAbd-xtcdFb .wvGCSb-F9IAbd-xtcdFb-LgbsSe.tk3N6e-LgbsSe.tk3N6e-LgbsSe { border-radius: 18px; height: auto; min-height: 36px; padding: 3px 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR { border-top: 1px solid rgb(232, 232, 232); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; padding: 18px 0px 7px; position: relative; outline: none; zoom: 1; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; padding: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-lCdvJf-fj0AZd { background-color: rgba(140, 196, 116, 0.5); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-gk6SMd-lCdvJf-fj0AZd { background-color: rgb(140, 196, 116); }

.HB1eCd-UMrnmb.HB1eCd-Guievd-WqyaDf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-lCdvJf-fj0AZd { background-color: highlight; color: highlighttext; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-dhWRR { border: 1px solid rgb(218, 220, 224); border-radius: 8px; margin: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR { border: 2px solid rgb(241, 243, 244); box-sizing: border-box; padding: 0px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .dhWRR-di8rgd-tJHJj.wvGCSb-dhWRR { border: 1px solid rgb(218, 220, 224); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-dhWRR:hover { background-color: rgb(254, 247, 224); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR:hover { background-color: transparent; border: 2px solid rgb(254, 239, 195); box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .dhWRR-di8rgd-tJHJj.wvGCSb-dhWRR:hover { border: 1px solid transparent; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YLEF4c { left: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YLEF4c { left: 0px; margin-top: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-SQuiCb .wvGCSb-W3vEtb-n0tgWb { position: absolute; top: 0px; right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-W3vEtb-n0tgWb > .wvGCSb-CTWaPd-j4gsHd { background-color: transparent; opacity: 0.7; }

.wvGCSb:not(.HB1eCd-UMrnmb).wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR:last-child { padding-bottom: 0px; }

.wvGCSb:not(.HB1eCd-UMrnmb).wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR:last-child .wvGCSb-dhWRR-nK2kYb { padding-bottom: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-pnL5fc-C58Yv { min-height: 48px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d { margin-right: 12px; min-height: 51px; padding: 0px 6px; position: relative; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-nhQw3d { margin-right: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d { margin-bottom: 8px; padding: 0px; top: 0px; }

.wvGCSb:not(.HB1eCd-UMrnmb).wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-nhQw3d { background-color: rgb(246, 246, 246); }

.wvGCSb:not(.HB1eCd-UMrnmb).wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-nhQw3d { background-color: rgb(255, 251, 225); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .HB1eCd-UMrnmb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe { background-color: rgb(241, 243, 244); border: 1px solid transparent; box-shadow: none; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover { background-color: rgb(241, 243, 244); box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .HB1eCd-UMrnmb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover { background-color: rgb(241, 243, 244); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover { border: 1px solid rgb(241, 243, 244); box-shadow: none; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd { background-color: rgb(241, 243, 244); box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb.HB1eCd-UMrnmb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd { background-color: rgb(241, 243, 244); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd { border: 1px solid rgb(232, 234, 237); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd { background-color: rgb(255, 251, 225); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd-bYHpTb { background-color: rgb(232, 240, 254); }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb.HB1eCd-UMrnmb .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd { background-color: rgb(254, 239, 195); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd { background-color: transparent; border: 2px solid rgb(253, 214, 99); box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; }

.wvGCSb.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .dhWRR-di8rgd-tJHJj.wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd { border: 1px solid transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc { margin-left: 60px; position: relative; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc { margin-left: 40px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc { margin-left: 0px; padding: 15px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od-biJjHb { -webkit-box-align: start; align-items: start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex-grow: 1; -webkit-box-pack: center; justify-content: center; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od-biJjHb .wvGCSb-dhWRR-oQLbGe { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 18px; letter-spacing: 0.25px; line-height: 20px; margin: 0px; max-width: 80%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-dhWRR-gqY2Od-biJjHb .wvGCSb-dhWRR-oQLbGe { max-width: 70%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od-biJjHb .wvGCSb-dhWRR-biJjHb { -webkit-box-align: center; align-items: center; color: rgb(95, 99, 104); display: flex; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 400; line-height: 16px; letter-spacing: 0.3px; margin: 0px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od-biJjHb > * { overflow: hidden; text-overflow: ellipsis; align-self: stretch; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-nhQw3d .wvGCSb-eKrold-TJEFFc { padding-top: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od { font-weight: 500; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .QpLw9-qnnXGd-lI7fHe .wvGCSb-dhWRR-gqY2Od { -webkit-box-align: center; align-items: center; display: inline-flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-RmniWd-mQXP { -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-align: center; align-items: center; background-color: rgb(26, 115, 232); border-radius: 9px; color: white; height: 16px; -webkit-box-pack: center; justify-content: center; margin: auto 0px; overflow: hidden; transform-origin: left center; transition: transform 0.2s ease-out 0s, color 0.1s ease-in 0s, border-radius 0.2s ease 0s, -webkit-transform 0.2s ease-out 0s; line-height: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-RmniWd-mQXP { margin-left: 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR:not(:hover) .wvGCSb-RmniWd-mQXP { border-radius: 50%; color: white; transform: scale(0.375); width: 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-gqY2Od span + .wvGCSb-RmniWd-mQXP { margin-left: 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR:not(:hover) .wvGCSb-RmniWd-Ne3sFf { color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-qJTHM { color: rgb(51, 51, 51); overflow-wrap: break-word; top: -7px; zoom: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-eKrold-qJTHM-haAclf { padding-top: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-biJjHb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-RDNXzf-Xhs9z { color: rgb(95, 99, 104); font-size: 12px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-biJjHb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-qrmfqe-bMcfAe { right: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-ZGNLv { color: rgb(204, 204, 204); font-size: 12px; line-height: 100%; padding: 0px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-nK2kYb { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; padding: 4px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-biJjHb:hover { text-decoration: underline; cursor: pointer; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-biJjHb:hover { text-decoration: none; cursor: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc { padding-right: 6px; margin-left: 30px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc { margin-left: 40px; padding-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-wTehdb-ORHb-haAclf { margin-left: -40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { background-color: rgb(255, 255, 255); border: 1px solid rgb(201, 212, 236); height: 23px; font-size: 12px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(60, 64, 67); font-size: 14px; line-height: 20px; min-height: 36px; padding: 8px; height: unset; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od:focus { border: 2px solid rgb(26, 115, 232); box-shadow: none; padding: 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-YPqjbf-BeDmAc.wvGCSb-YPqjbf-YsTx5 .wvGCSb-YPqjbf-B7I4Od { background-color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-DyVDA-BeDmAc .wvGCSb-YPqjbf-B7I4Od { height: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-MGbz6c { margin: 4px 12px 3px 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-MGbz6c { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d { background-color: rgb(239, 242, 249); border-radius: 0px 0px 6px 6px; padding: 6px 0px 2px 6px; position: relative; zoom: 1; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d { background-color: white; border: 1px solid rgb(218, 220, 224); border-radius: 4px; padding: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d { background: inherit; border: 1px solid transparent; margin: 0px; padding: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-dhWRR-xuvf2d { background: inherit; border: 1px solid transparent; left: -40px; margin: 0px; padding: 0px; width: 110%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-xuvf2d { background-color: rgb(246, 246, 246); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-xuvf2d { background-color: white; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-xuvf2d { background: inherit; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-xuvf2d { background: inherit; left: -40px; width: 110%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-xuvf2d { left: 0px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-MZArnb { position: absolute; right: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-MZArnb .wvGCSb-no16zc-ldDtVd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-MZArnb .wvGCSb-ERydpb-ldDtVd { height: 28px; margin: 0px; position: relative; top: auto; right: auto; display: inline-block; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-MZArnb { right: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe .wvGCSb-dhWRR-MZArnb { right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-KjQ5hb-n0tgWb { position: absolute; right: -12px; top: 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-qrmfqe-bMcfAe { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-qrmfqe-bMcfAe > .wvGCSb-pnL5fc-qrmfqe { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 12px; font-weight: 500; color: rgb(17, 85, 204); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-jNm5if-bMcfAe > .wvGCSb-pnL5fc-jNm5if, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-WlKKfd-bMcfAe > .wvGCSb-pnL5fc-WlKKfd { color: rgb(153, 153, 153); line-height: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-jNm5if-bMcfAe > .wvGCSb-pnL5fc-jNm5if:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-qrmfqe-bMcfAe > .wvGCSb-pnL5fc-qrmfqe:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-WlKKfd-bMcfAe > .wvGCSb-pnL5fc-WlKKfd:hover { text-decoration: underline; cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d:hover .wvGCSb-pnL5fc-jNm5if, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d:hover .wvGCSb-pnL5fc-WlKKfd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-pnL5fc-jNm5if, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-pnL5fc-WlKKfd { color: rgb(17, 85, 204); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(241, 243, 244); border-top-left-radius: 8px; border-top-right-radius: 8px; margin: -1px; outline: none; padding: 10px 16px; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR:hover .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(254, 239, 195); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(253, 214, 99); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR:hover .wvGCSb-dhWRR-tJHJj-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd.wvGCSb-dhWRR .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(218, 220, 224); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-haAclf { display: inline-flex; min-width: 0px; -webkit-box-flex: 1; flex: 1 1 0%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-dwJgKd-T3yXSc { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-dwJgKd-P86uke { color: rgb(60, 64, 67); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-auswjd .dhWRR-tJHJj-dwJgKd-P86uke { color: rgb(32, 33, 36); font-weight: bold; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-dwJgKd-tJHJj, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-auswjd .dhWRR-tJHJj-T3yXSc-KoToPc .dhWRR-tJHJj-dwJgKd-T3yXSc { display: block; width: 90%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj { display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-EvNWZc .dhWRR-tJHJj { width: 90%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-auswjd .dhWRR-tJHJj-T3yXSc-KoToPc .dhWRR-tJHJj { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-auswjd .dhWRR-tJHJj-T3yXSc-KoToPc .dhWRR-tJHJj div { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-pnL5fc-auswjd .dhWRR-tJHJj-T3yXSc-KoToPc .dhWRR-tJHJj .dhWRR-tJHJj-P86uke { overflow: hidden; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-KoToPc .dhWRR-tJHJj .dhWRR-tJHJj-T3yXSc { overflow-wrap: break-word; white-space: normal; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-clz4Ic-haAclf { display: inline-flex; -webkit-box-align: center; align-items: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-clz4Ic-haAclf .dhWRR-tJHJj-clz4Ic { padding: 0px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-P86uke-haAclf { -webkit-box-align: center; align-items: center; display: inline-flex; font-weight: 500; min-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-P86uke-haAclf.tJHJj-SfQLQb-T3yXSc { max-width: 50%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj .dhWRR-tJHJj-T3yXSc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-P86uke-haAclf .dhWRR-tJHJj-qdIk2c-P86uke { line-height: 20px; max-height: 20px; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-P86uke-haAclf .dhWRR-tJHJj-qdIk2c-clz4Ic { margin-right: 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-c6xFrd-haAclf { cursor: pointer; display: none; position: absolute; right: 0px; top: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-EvNWZc .dhWRR-tJHJj-T3yXSc-c6xFrd-haAclf { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-EvNWZc .dhWRR-tJHJj-T3yXSc-vhaaFf-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-KoToPc.dhWRR-tJHJj-EvNWZc .dhWRR-tJHJj-T3yXSc-KoToPc-LgbsSe { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-KoToPc.dhWRR-tJHJj-EvNWZc .dhWRR-tJHJj-T3yXSc-vhaaFf-LgbsSe { display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR { border-radius: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-dhWRR { border: none; outline: rgb(199, 199, 199) solid 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb.wvGCSb-F6aDIf .wvGCSb-dhWRR:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover { border: none; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 2px, rgba(0, 0, 0, 0.15) 0px 2px 6px 2px; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb.wvGCSb.wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd { border: none; box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd { background-color: rgb(242, 242, 242); box-shadow: rgba(0, 0, 0, 0.3) 0px 1px 3px, rgba(0, 0, 0, 0.15) 0px 4px 8px 3px; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .dhWRR-tJHJj, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .dhWRR-tJHJj-dwJgKd-P86uke, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf .wvGCSb-gkA7Yd-Wz3zdc-T3yXSc-cHYyed { font: 500 12px / 16px "Google Sans", Roboto, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-tJHJj-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background: rgb(242, 242, 242); border-top-left-radius: 11px; border-top-right-radius: 11px; margin: 0px; padding: 6px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR:hover .wvGCSb-dhWRR-tJHJj-haAclf { background: rgb(255, 240, 209); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-dhWRR-tJHJj-haAclf { background: rgb(255, 187, 41); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover { background: rgb(242, 242, 242); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR:hover .wvGCSb-dhWRR-tJHJj-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd.wvGCSb-dhWRR .wvGCSb-dhWRR-tJHJj-haAclf { background-color: rgb(227, 227, 227); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb .wvGCSb-dhWRR-bN97Pc { padding: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId { border-radius: 11px 11px 0px 0px; margin: 1px; padding: 10px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .wvGCSb-dhWRR-tJHJj-haAclf + .wvGCSb-dhWRR-bN97Pc .wvGCSb-GpPaId { border-radius: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-MZArnb { opacity: 0; transition: opacity 0.25s cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-MZArnb { opacity: 0; transition: opacity 0.25s cubic-bezier(0.4, 0, 0.2, 1) 0s; -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-MZArnb div[role="button"] { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-W3vEtb-n0tgWb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR-MZArnb:focus-within, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR:hover .wvGCSb-dhWRR-MZArnb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR:focus .wvGCSb-dhWRR-MZArnb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-dhWRR-MZArnb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR:hover .wvGCSb-gkA7Yd-Wz3zdc-MZArnb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR:focus .wvGCSb-gkA7Yd-Wz3zdc-MZArnb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-MZArnb { opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .HB1eCd-UMrnmb .wvGCSb-dhWRR-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { border-radius: 18px; padding: 8px 7px 8px 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-F6aDIf .dhWRR-tJHJj-T3yXSc-c6xFrd-haAclf { top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .dhWRR-tJHJj-T3yXSc-c6xFrd-haAclf .HB1eCd-HzV7m-LgbsSe { border-radius: 100%; display: flex; height: 32px; -webkit-box-pack: center; justify-content: center; width: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-gkA7Yd-Wz3zdc-haAclf { display: flex; -webkit-box-align: center; align-items: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-oQLbGe { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-bN97Pc .wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-oQLbGe .wvGCSb-oQLbGe { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 18px; letter-spacing: 0.25px; line-height: 20px; margin: 0px; max-width: 80%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-Wz3zdc { height: 18px; width: 18px; margin-right: 10px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-xtcdFb-Wz3zdc.wvGCSb-gkA7Yd-Wz3zdc-Wz3zdc-sLO9V-qnnXGd { font-family: "Noto Color Emoji", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 17px; margin-top: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-bN97Pc { padding-left: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-tL9eOd { display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-Wz3zdc-nUpftc-YLEF4c { left: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf .wvGCSb-gkA7Yd-Wz3zdc-T3yXSc-cHYyed { line-height: 20px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-style: normal; font-size: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(241, 243, 244); display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-align: center; align-items: center; padding: 10px 16px; border-top-left-radius: 8px; border-top-right-radius: 9px; margin: -1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc-JIbuQc-haAclf { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; position: relative; padding-bottom: 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-FDWhSe { color: rgb(128, 134, 139); font-size: 11px; font-style: italic; text-align: left; white-space: pre-wrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .gkA7Yd-Wz3zdc-lI7fHe-nUpftc-tJHJj-clz4Ic { padding: 0px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :not(docos-docoview-resolved) .wvGCSb-dhWRR:hover .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(254, 239, 195); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb :not(docos-docoview-resolved) .wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(253, 214, 99); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR.wvGCSb-pnL5fc-IIEkAe:hover .wvGCSb-gkA7Yd-Wz3zdc-tJHJj-haAclf { background-color: rgb(218, 220, 224); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR.wvGCSb-pnL5fc-auswjd .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc { background-color: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-MZArnb { position: absolute; right: 0px; top: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { margin: 0px 8px 0px 0px; width: 28px; height: 28px; vertical-align: middle; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-W3vEtb-n0tgWb .VIpgJd-INgbqf-xl07Ob-LgbsSe-n0tgWb-Q4BLdf { min-width: 14px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-gkA7Yd-Wz3zdc-lI7fHe-nUpftc-j4LONd-cnfHN { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 18px; letter-spacing: 0.25px; line-height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-gkA7Yd-Wz3zdc-MZArnb { display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-pack: center; justify-content: center; background: none; border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background: none rgba(68, 71, 70, 0.08); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf .wvGCSb-dhWRR .wvGCSb-gkA7Yd-Wz3zdc-WlKKfd-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background: none rgba(68, 71, 70, 0.12); border-radius: 100%; height: 32px; width: 32px; border: 1px solid transparent !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue .wvGCSb-YPqjbf-LgbsSe-oKdM2c { padding-bottom: 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue .wvGCSb-YPqjbf-aIWppb { margin: 0px 4px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue .wvGCSb-YPqjbf-IbE0S { background: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-PvRhvb-Bz112c { display: flex; -webkit-box-align: center; align-items: center; margin-right: 12px; height: 24px; width: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-PvRhvb-Bz112c .HB1eCd-UMrnmb-PvRhvb-Bz112c-r9oPif { height: 24px; margin: 0px; width: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-PvRhvb-Bz112c-Jt5cK { fill: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-haAclf { line-height: 140%; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-bN97Pc { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-PLt2Ue-bN97Pc { position: static; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-XHP5j { color: rgb(17, 85, 204); cursor: pointer; font-size: 12px; position: absolute; right: 0px; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-XHP5j:hover { text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PrY1nf .wvGCSb-PLt2Ue-XHP5j { color: rgb(153, 153, 153); cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PrY1nf .wvGCSb-PLt2Ue-XHP5j:hover { text-decoration: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-QCAl5e { bottom: -10px; color: rgb(17, 85, 204); cursor: pointer; font-size: 12px; padding-right: 5px; padding-top: 5px; position: absolute; right: 5px; text-decoration: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PrY1nf .wvGCSb-PLt2Ue-QCAl5e { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-I1HBjd { color: rgb(51, 51, 51); padding: 12px 0px 12px 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-cD65uc { background-color: rgb(254, 247, 224); border-top: 1px solid rgb(218, 220, 224); border-bottom: 1px solid rgb(218, 220, 224); color: rgb(95, 99, 104); font-weight: 500; padding: 12px 20px; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-Q5sUsf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-Q5sUsf:visited { color: rgb(26, 115, 232); font-weight: 400; margin-left: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-cD65uc { border-top: 0px; box-sizing: border-box; height: 62px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-SvJh7b { margin: 6px 29px 10px 20px; position: relative; zoom: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-SvJh7b-bN97Pc { margin-left: 61px; position: relative; zoom: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xqKM5b { font-size: 12px; font-weight: 500; margin-bottom: 3px; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-r4nke { font-size: 1.2em; margin: 20px 5px 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-YPqjbf-BeDmAc { top: -4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-YPqjbf-BeDmAc .wvGCSb-YPqjbf-aIWppb { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-YPqjbf-BeDmAc .wvGCSb-YPqjbf-B7I4Od { font-size: 12px; height: 30px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-WS1epc-xtcdFb-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-eMXQ4e-F8G5oc-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-lQVAed-Ne3sFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-xuvf2d .wvGCSb-YPqjbf-TJEFFc-Ne3sFf { color: rgb(119, 119, 119); line-height: normal; margin-top: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-u0pjoe { background-color: rgb(221, 75, 57); border: 1px solid rgb(96, 32, 25); border-radius: 4px; color: rgb(255, 255, 255); margin: 6px; padding: 6px; text-align: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj { -webkit-box-align: center; align-items: center; display: flex; background-color: rgb(245, 245, 245); max-height: 52px; overflow: hidden; padding: 10px 29px 10px 20px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj { background-color: white; border-bottom: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj-I5GmGe-ma6Yeb-vFHz9d { border-radius: 8px 8px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .HB1eCd-UMrnmb .wvGCSb-PLt2Ue-tJHJj { padding: 12px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe { margin-right: 4px; width: 40px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe { border-radius: 50%; height: 40px; margin: 0px; padding: 4px; width: 40px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe.HB1eCd-HzV7m-LgbsSe-XpnDCe { line-height: 32px; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-ZmdkE.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-XpnDCe.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GUUVJe-EnFNjd-LgbsSe .HB1eCd-HzV7m-LgbsSe-auswjd.HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae { background-color: rgb(232, 234, 237); border: none; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-LgbsSe .HB1eCd-HzV7m-LgbsSe-bN97Pc { top: 5px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { -webkit-box-align: center; align-items: center; border-radius: 50%; display: flex; height: 32px; -webkit-box-pack: center; justify-content: center; margin: 0px; min-width: 32px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { padding: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { display: inline-block; float: left; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-jNm5if-r4nke-haAclf { -webkit-box-align: center; align-items: center; display: flex; margin-right: auto; order: -1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-F6aDIf .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS.wvGCSb-jNm5if-tJHJj-r4nke { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 16px; font-weight: 500; line-height: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .wvGCSb-yOOK0-EnFNjd { padding: 0px 0px 0px 10px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-PLt2Ue-tJHJj .wvGCSb-yOOK0-EnFNjd { padding: 0px; width: 160px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe { border-color: transparent; background-color: transparent; background-image: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-auswjd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-XpnDCe { border-color: rgb(198, 198, 198); background-color: rgb(248, 248, 248); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(248, 248, 248)), to(rgb(241, 241, 241))); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { visibility: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-auswjd .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { visibility: visible; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .wvGCSb-GmVRCe-cHYyed-Bz112c { opacity: 0.3; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GmVRCe-cHYyed { -webkit-box-align: center; align-items: center; display: flex; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-Bz112c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-GmVRCe-cHYyed-Bz112c { margin: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-tJHJj .tk3N6e-LgbsSe-OWB6Me .wvGCSb-RmniWd-jNm5if-Bz112c { opacity: 0.15; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-haAclf { -webkit-box-align: center; align-items: center; border-bottom: 1px solid rgb(218, 220, 224); box-sizing: border-box; display: none; -webkit-box-pack: justify; justify-content: space-between; max-height: 0px; overflow: hidden; padding: 0px 20px; transition: max-height 0.3s ease-in-out 0s, padding 0.3s ease-in-out 0s; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-FNFY6c { display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-PBWx0c { max-height: 100px; padding: 10px 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe { width: 75%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe .wvGCSb-PLt2Ue-G0jgYd-YPqjbf { border: 1px solid rgb(189, 193, 198); border-radius: 8px; box-sizing: border-box; height: auto; padding: 8px 10px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe .wvGCSb-PLt2Ue-G0jgYd-YPqjbf:focus { border-color: rgb(77, 144, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe { margin-right: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe .HB1eCd-HzV7m-LgbsSe-Kb3HCc-zTETae.HB1eCd-HzV7m-LgbsSe-ZmdkE { background-color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-LgbsSe .HB1eCd-HzV7m-LgbsSe-ksKsZd-PQbLGe { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-xxlfEe-TvD9Pc-Bz112c-SxQuSe { width: 18px; height: 18px; margin: 1px 2px 2px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Bz112c.HB1eCd-HzV7m.wvGCSb-PLt2Ue-GUUVJe-EnFNjd-Bz112c-SxQuSe { width: 24px; height: 24px; margin: 1px 2px 2px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RXQi4b-HB1eCd-tJHJj .wvGCSb-gkA7Yd-nUpftc { position: relative; overflow: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RXQi4b-HB1eCd-tJHJj .wvGCSb-gkA7Yd-nUpftc-NBtyUd { max-height: 369px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RXQi4b-HB1eCd-tJHJj:not(.HB1eCd-UMrnmb) .wvGCSb-gkA7Yd-nUpftc > .wvGCSb-dhWRR:first-child { border-top-color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-gkA7Yd-nUpftc { bottom: 1px; max-height: none; overflow: hidden auto; position: absolute; top: 116px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-iQd6Fc.wvGCSb-gkA7Yd-nUpftc { margin-top: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb-bN97Pc .wvGCSb-gkA7Yd-nUpftc.s4YTVd-NBtyUd-IT5dJd-ORHb { top: 170px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-Bz112c { display: inline-block; vertical-align: middle; margin: 4px 5px 5px 2px; opacity: 0.65; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-Bz112c { opacity: 1; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe { box-shadow: none; background-color: white; background-image: none; cursor: pointer; border-radius: 2px; border-width: initial; border-style: none; border-image: initial; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 500; line-height: 16px; padding: 2px 6px 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe { background-color: transparent; color: transparent; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { border-radius: 50%; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { box-shadow: none; background-color: rgb(232, 240, 254); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-ZmdkE { background-color: rgb(241, 243, 244); border-radius: 50%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-XpnDCe { background-color: rgb(232, 234, 237); border-radius: 50%; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd { box-shadow: none; background-color: rgb(210, 227, 252); background-image: none; cursor: pointer; border-radius: 2px; border-width: 1px; border-color: transparent !important; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-auswjd { background-color: rgb(232, 234, 237); outline: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { font-family: "Google Sans"; font-size: 14px; font-weight: 500; line-height: 28px; text-transform: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { -webkit-box-align: center; align-items: center; color: rgb(60, 64, 67); font-family: "Google Sans"; font-size: 14px; font-weight: 500; line-height: 28px; text-transform: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { -webkit-box-align: center; align-items: center; border: 1px solid rgb(218, 220, 224); border-radius: 24px; color: rgb(95, 99, 104); display: flex; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf { background-color: rgb(232, 240, 254); border: none; color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.HB1eCd-UMrnmb.HB1eCd-v3pZbf-yQ1rOb-Bz112c-n9v5ye.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c-RJLb9c { filter: brightness(0) saturate(100%) invert(28%) sepia(99%) saturate(2090%) hue-rotate(205deg) brightness(98%) contrast(86%); content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_gm3_grey_medium.svg"); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae.yOOK0-x9Ufpf .HB1eCd-Bz112c { display: inline-block; margin-bottom: 4px; margin-right: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae .HB1eCd-Bz112c { display: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-cHYyed { margin-left: 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-cHYyed { overflow: hidden; text-overflow: ellipsis; white-space: nowrap; width: 100px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { color: rgb(32, 33, 36); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { color: rgb(24, 90, 188); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { color: rgb(24, 90, 188); background-color: rgb(248, 251, 255); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { background-color: rgb(233, 241, 254); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd { background-color: rgb(225, 236, 254); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE { background: rgba(60, 64, 67, 0.04); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { background: rgba(60, 64, 67, 0.12); border: 1px solid rgb(32, 33, 36); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd { background: rgba(60, 64, 67, 0.16); border: 1px solid rgb(218, 220, 224); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(95, 99, 104); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(32, 33, 36); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-auswjd .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd .yOOK0-x9Ufpf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-ZmdkE .HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-j4gsHd-Bz112c { fill: rgb(24, 90, 188); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd-Guievd-WqyaDf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae-XpnDCe { filter: invert(100%); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-yOOK0-EnFNjd-Guievd-WqyaDf.HB1eCd-HzV7m-xl07Ob-LgbsSe-Kb3HCc-zTETae { outline: transparent solid 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-bN97Pc .wvGCSb-jNm5if-fmcmS { padding: 2px 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-LgbsSe.tk3N6e-LgbsSe-OWB6Me { background-color: white; color: rgb(241, 243, 244); cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld { cursor: grab; border-color: rgb(232, 234, 237); border-style: solid; border-width: 1px 0px 0px; height: 8px; width: 100%; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld-Bz112c { height: 4px; margin: 2px auto 0px; width: 20px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-haAclf .PLt2Ue-CCJ0ld:hover { background-color: rgb(232, 234, 237); cursor: grab; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-NkyfNe-imnzkf-m9bMae-MJoBVe-bN97Pc { color: rgb(128, 134, 139); padding-top: 24px; text-align: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-Bz112c { display: inline-block; vertical-align: middle; margin: 4px 5px 5px 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-Bz112c { margin-left: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-UMrnmb-b3rLgd-Bz112c-Jt5cK, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-Bz112c-Jt5cK { fill: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-UMrnmb-b3rLgd-Bz112c-Jt5cK, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-G0jgYd-RDNXzf-Bz112c-Jt5cK, .HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-RmniWd-jNm5if-Bz112c-Jt5cK, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-UMrnmb-b3rLgd-Bz112c-Jt5cK, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-G0jgYd-RDNXzf-Bz112c-Jt5cK, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-RmniWd-jNm5if-Bz112c-Jt5cK { fill: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-OWB6Me .wvGCSb-RmniWd-jNm5if-Bz112c-Jt5cK { fill: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed { text-align: left; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed { height: 27px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-fmcmS { display: inline-block; height: 17px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-fmcmS { line-height: 16px; height: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-GmVRCe-cHYyed-LwH6nd { visibility: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe { -webkit-box-align: center; align-items: center; background-color: rgb(255, 255, 255); bottom: 1px; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; -webkit-box-pack: justify; justify-content: space-between; max-height: none; position: absolute; text-align: center; top: 116px; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-tJHJj-HiaYvf { height: 200px; margin-top: 2vh; width: 300px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-bN97Pc-htvI8d-jNm5if { margin-bottom: 16px; color: rgb(60, 64, 67); font-size: 14px; font-weight: 400; letter-spacing: 0.2px; line-height: 20px; width: 158px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-htvI8d-jNm5if-LgbsSe.HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe { text-transform: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-yePe5c { letter-spacing: 0.2px; font-size: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-yePe5c-D1hqkb { color: rgb(128, 134, 139); font-weight: 500; line-height: 18px; margin-bottom: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-PLt2Ue-x5ghY-MJoBVe-yePe5c-D1hqkb-WjNrPc { color: rgb(128, 134, 139); font-weight: 400; font-size: 12px; line-height: 18px; width: 191px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb { background-color: rgb(239, 242, 249); color: rgb(102, 102, 102); font-size: 12px; padding: 6px 6px 0px; position: relative; margin-bottom: 3px; min-height: 24px; outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d { outline: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb { background-color: white; border: 1px solid rgb(218, 220, 224); border-radius: 4px; font-size: 14px; margin-bottom: 8px; padding: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb { background: inherit; border: 1px solid transparent; margin: 0px; padding: 8px 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-SQuiCb { background: inherit; border: 1px solid transparent; left: -40px; margin: 0px; padding: 8px 0px; width: 110%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb { left: 0px; width: 100%; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d-bN97Pc { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-SQuiCb { background-color: rgb(246, 246, 246); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-SQuiCb { background-color: white; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-SQuiCb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-pnL5fc-IIEkAe .wvGCSb-SQuiCb { background: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-YLEF4c { left: 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-YLEF4c { left: 16px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-YLEF4c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-SQuiCb-YLEF4c { left: 0px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d-bN97Pc { padding-left: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-bN97Pc { padding-left: 30px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-bN97Pc { padding-left: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-oQLbGe { color: black; font-weight: 500; }

.wvGCSb:not(.HB1eCd-UMrnmb).wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-oQLbGe { left: -2px; margin: 0px 4px; right: -2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .QpLw9-qnnXGd-lI7fHe .wvGCSb-SQuiCb-oQLbGe { -webkit-box-align: center; align-items: center; display: inline-flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-oQLbGe { color: rgb(60, 64, 67); letter-spacing: 0.25px; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; line-height: 20px; padding-right: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb .wvGCSb-RmniWd-mQXP { -webkit-box-flex: 0; flex: 0 0 auto; -webkit-box-align: center; align-items: center; background-color: rgb(26, 115, 232); border-radius: 9px; color: white; height: 16px; -webkit-box-pack: center; justify-content: center; margin: auto 0px; overflow: hidden; transform-origin: left center; transition: transform 0.2s ease-out 0s, color 0.1s ease-in 0s, border-radius 0.2s ease 0s, -webkit-transform 0.2s ease-out 0s; line-height: 16px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb:not(:hover) .wvGCSb-RmniWd-mQXP { border-radius: 50%; color: white; transform: scale(0.375); width: 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb span + .wvGCSb-RmniWd-mQXP { margin-left: 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb:not(:hover) .wvGCSb-RmniWd-Ne3sFf { color: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-qJTHM { color: rgb(51, 51, 51); margin: 0px; top: -4px; width: 100%; overflow-wrap: break-word; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-fmcmS, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-biJjHb { position: relative; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-fmcmS { width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-FDWhSe { padding-bottom: 4px; font-style: italic; color: rgb(153, 153, 153); font-size: 11px; white-space: pre; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-biJjHb { color: rgb(153, 153, 153); font-size: 11px; white-space: pre; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-FDWhSe.wvGCSb-SQuiCb-FDWhSe { white-space: pre-wrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-SQuiCb .wvGCSb-eKrold-bMcfAe { display: inline; top: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-DyVDA-BeDmAc .wvGCSb-YPqjbf-B7I4Od { height: 23px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-eKrold-T3yXSc { border-left: 1px solid rgb(204, 204, 204); font-style: italic; font-size: 12px; padding: 3px 10px; position: relative; zoom: 1; overflow-wrap: break-word; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR .wvGCSb-eKrold-T3yXSc { margin: 8px 0px; padding: 0px 8px 0px 16px; border-left-width: 3px; border-left-color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-cHYyed { font-size: 11px; font-weight: 500; color: rgb(153, 153, 153); margin-right: 2px; padding: 0px; }

.HB1eCd-UMrnmb.wvGCSb-F6aDIf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb-YLEF4c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-wvGCSb-Z0Arqf-PvRhvb .wvGCSb-SQuiCb-YLEF4c { font-size: 12px; overflow-wrap: break-word; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-cHYyed { color: rgb(60, 64, 67); letter-spacing: 0.8px; line-height: 21px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; text-transform: uppercase; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-qAWA2 { overflow: hidden; height: 18px; padding-left: 3px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-vhaaFf { height: 21px; padding-left: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-KoToPc { background: rgb(255, 255, 255); padding: 3px 5px 0px; position: absolute; right: 0px; top: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-KoToPc { padding: 0px 5px 0px 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-vhaaFf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-KoToPc { color: rgb(17, 85, 204); visibility: hidden; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-vhaaFf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-KoToPc { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-T3yXSc-vhaaFf { visibility: visible; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd .wvGCSb-eKrold-T3yXSc-KoToPc { visibility: visible; background: rgb(255, 251, 225); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-vhaaFf:hover, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-eKrold-T3yXSc-KoToPc:hover { cursor: pointer; text-decoration: underline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d .wvGCSb-JIbuQc-fmcmS, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb .wvGCSb-JIbuQc-fmcmS { color: rgb(119, 119, 119); font-style: italic; overflow-wrap: break-word; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d .wvGCSb-JIbuQc-fmcmS, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-SQuiCb .wvGCSb-JIbuQc-fmcmS { color: rgb(60, 64, 67); opacity: 0.7; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-nhQw3d .wvGCSb-JIbuQc-fmcmS { display: inline-block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-dhWRR-bN97Pc .wvGCSb-YPqjbf-lQVAed-b0t70b { margin-top: -5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b { -webkit-box-align: center; align-items: center; border-radius: 8px; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; padding: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-Tswv1b { background: rgb(232, 240, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-Tswv1b > .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_blue.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-lHjamb { background: rgb(254, 239, 195); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-GMvhG { background: rgb(251, 188, 4); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-lHjamb > .HB1eCd-Bz112c-RJLb9c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-GMvhG > .HB1eCd-Bz112c-RJLb9c { content: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_dark.svg"); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b > .HB1eCd-Bz112c { flex-shrink: 0; height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Hn6s1b-Ne3sFf { color: rgb(32, 33, 36); font: 400 14px / 20px Roboto, sans-serif; letter-spacing: 0.2px; margin-left: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-suEOdc { display: inline-block; max-width: 35ch; text-align: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc { box-sizing: border-box; text-align: left; width: 330px; }

.wvGCSb-XS83If-bN97Pc.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb { border-radius: 8px; white-space: normal; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc .HB1eCd-Hn6s1b { margin-bottom: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc [role="heading"] { color: rgb(32, 33, 36); font: 400 18px / 24px "Google Sans", sans-serif; margin-bottom: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc p { color: rgb(95, 99, 104); font: 500 11px / 16px Roboto, sans-serif; letter-spacing: 0.8px; margin-bottom: 16px; text-transform: uppercase; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf { padding: 0px; display: block; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf.tk3N6e-Ru3Ixf-OWB6Me { opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf + .tk3N6e-Ru3Ixf { margin-top: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-GCYh9b { border: 2px solid rgb(95, 99, 104); height: 15px; width: 15px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-GCYh9b { left: 3px; top: 50%; transform: translateY(-50%) scale(1.2); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-ZmdkE:not(.tk3N6e-Ru3Ixf-OWB6Me) .tk3N6e-Ru3Ixf-GCYh9b { cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-GCYh9b::before { border-color: transparent; border-radius: 50%; border-style: solid; border-width: 6px; content: ""; height: 19px; left: -10.5px; position: absolute; top: -10.5px; transform: scale(0.8333); width: 19px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc :not(.tk3N6e-Ru3Ixf-OWB6Me):not(.tk3N6e-Ru3Ixf-XpnDCe) .tk3N6e-Ru3Ixf-GCYh9b:hover::before { border-color: rgba(0, 0, 0, 0.06); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-XpnDCe .tk3N6e-Ru3Ixf-GCYh9b::before { border-color: rgb(232, 240, 254); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie .tk3N6e-Ru3Ixf-GCYh9b { border-color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie.tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-GCYh9b::after { background-color: rgb(26, 115, 232); border-color: rgb(26, 115, 232); border-width: 2px; height: 7px; left: 2px; margin: 0px; top: 2px; width: 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf .tk3N6e-Ru3Ixf-V67aGc { margin-left: 36px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-V67aGc label { color: rgb(60, 64, 67); display: block; font: 500 14px / 24px "Google Sans", sans-serif; letter-spacing: 0.1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-barxie .tk3N6e-Ru3Ixf-V67aGc label { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-GCYh9b-LgbsSe-JNdkSc .tk3N6e-Ru3Ixf-V67aGc span { color: rgb(95, 99, 104); font: 400 12px / 16px Roboto, sans-serif; letter-spacing: 0.3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-XS83If-bN97Pc hr { border-right: none; border-bottom: none; border-left: none; border-image: initial; border-top: 1px solid rgb(189, 193, 198); margin: 16px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-B7I4Od { margin: 0px; padding: 2px; font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; resize: none; outline-width: 0px !important; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Jiyx5 { list-style: none; margin: 0px; padding: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Jiyx5:focus { outline: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL { background: rgb(255, 255, 255); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .MsdWL { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.nhiZfc { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; height: 48px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.nhiZfc .E8WqE { height: 24px; width: 24px; margin-right: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.XdSAtd { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; height: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.XdSAtd .E8WqE { height: 20px; width: 20px; margin-right: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.HddOwd { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; height: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.HddOwd .E8WqE { height: 20px; width: 20px; margin-right: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL:hover { background: rgba(10, 10, 10, 0.04); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .MsdWL:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MsdWL.qs41qe { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .MsdWL.qs41qe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.25), rgba(232, 234, 237, 0.25)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .jcbibd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; max-width: 450px; padding-left: 12px; padding-right: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .w8bLS { -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .B92god { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hMC4ff { -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .E8WqE { margin-left: 0px; }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .E8WqE { filter: brightness(0) invert(1); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EKzqb { color: rgb(60, 64, 67); text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .EKzqb { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .bylmg { color: rgb(95, 99, 104); margin-left: 48px; margin-right: 0px; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .bylmg { color: rgb(218, 220, 224); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .heO6Yc { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 4px; outline: transparent solid 1px; overflow: hidden; padding-bottom: 8px; padding-top: 8px; position: absolute; user-select: none; z-index: 999999; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .heO6Yc .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .heO6Yc { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O5UuBc { font-family: "Google Sans", Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; color: rgb(26, 115, 232); -webkit-box-align: center; align-items: center; background: none; border-radius: 4px; border: none; outline: transparent solid 1px; display: flex; height: 36px; line-height: unset; padding: 0px 8px; user-select: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .O5UuBc { color: rgb(138, 180, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O5UuBc:hover { background-color: rgba(26, 115, 232, 0.04); color: rgb(23, 78, 166); cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .O5UuBc:hover { background-color: rgba(138, 180, 248, 0.04); color: rgb(210, 227, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O5UuBc:focus { background-color: rgba(26, 115, 232, 0.12); color: rgb(23, 78, 166); cursor: pointer; outline-width: 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .O5UuBc:focus { background-color: rgba(138, 180, 248, 0.12); color: rgb(210, 227, 252); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O5UuBc.RDPZE { color: rgba(60, 64, 67, 0.38); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .O5UuBc.RDPZE { color: rgba(232, 234, 237, 0.38); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O5UuBc.RDPZE:focus { background-color: rgba(60, 64, 67, 0.12); color: rgba(60, 64, 67, 0.38); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .O5UuBc.RDPZE:focus { background-color: rgba(232, 234, 237, 0.12); color: rgba(232, 234, 237, 0.38); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .q5Gute { -webkit-box-align: center; align-items: center; background: rgba(32, 33, 36, 0.6); box-sizing: border-box; display: flex; height: 100%; -webkit-box-pack: center; justify-content: center; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 999999; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .qnxR0c { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .qnxR0c { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .cySkyb { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 8px; max-width: 300px; outline: transparent solid 1px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .cySkyb .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .cySkyb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h6zUze { margin: 24px 24px 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tAzG6 { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .g9hvRc { width: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .xQiMxd { -webkit-box-align: center; align-items: center; background: rgba(32, 33, 36, 0.6); box-sizing: border-box; display: flex; height: 100%; -webkit-box-pack: center; justify-content: center; left: 0px; position: fixed; top: 0px; width: 100%; z-index: 999999; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .mSjfjb { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .mSjfjb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tFDhVb { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 500; color: rgb(32, 33, 36); margin: 24px 24px 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .tFDhVb { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EoolDb { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 8px; max-width: 300px; outline: transparent solid 1px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EoolDb .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .EoolDb { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Pmtn0b { margin: 24px 24px 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .X23yUb { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(60, 64, 67); margin-bottom: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .X23yUb { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ADqTKb { color: rgb(26, 115, 232); text-decoration: underline; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .ADqTKb { color: rgb(138, 180, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ADqTKb:visited { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .ADqTKb:visited { color: rgb(138, 180, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tlQjad { display: flex; -webkit-box-pack: end; justify-content: flex-end; padding: 8px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .mtq6kd { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .A6DTme { border-radius: 50%; outline: transparent solid 1px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hIJ6Le { margin: auto; display: block; height: 100%; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .vi1cfb { position: absolute; bottom: 0px; right: 0px; display: none; height: 30%; width: 30%; min-height: 30%; min-width: 30%; object-fit: cover; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .vi1cfb.ZiwkRe { display: inline; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .KKjvXb .vi1cfb { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .PS6m6 { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; height: inherit; width: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aGbmDb { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 0%; overflow: hidden; height: inherit; -webkit-box-align: stretch; align-items: stretch; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AcwQxb { display: flex; -webkit-box-flex: 1; flex: 1 1 0%; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IW1j2d { margin: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Khf4w { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-flex: 1; flex: 1 1 auto; -webkit-box-align: center; place-items: center; transition: background 50ms ease-in-out 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Khf4w.JpY6Fd { background-clip: padding-box; background-color: rgb(189, 193, 198); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ew7bve { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .k8rr2e .ew7bve { display: block; fill: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .k8rr2e .ew7bve { fill: rgb(154, 160, 166); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .ZlXryd { opacity: 1; display: block; transition: opacity 50ms ease-in-out 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .JpY6Fd .ZlXryd { opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .k8rr2e .ZlXryd { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AGaBze { background: rgb(255, 255, 255); border-bottom: 1px solid rgb(218, 220, 224); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AGaBze { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .haq1x { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; padding: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .rr5U0b { -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tJRcje { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XsnHSd { align-content: flex-start; -webkit-box-align: start; align-items: flex-start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-flow: column nowrap; margin-left: 12px; margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .RWXYif { -webkit-box-flex: initial; flex: initial; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .awj5uc { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; color: rgb(32, 33, 36); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .awj5uc { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .J7kVrb { font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; color: rgb(60, 64, 67); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .J7kVrb { color: rgb(154, 160, 166); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .fasgab { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .vG6Gfe { height: inherit; position: relative; width: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .L7D8v { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aAzAef { margin-bottom: 20px; font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .aAzAef { color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .TeNodb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; color: rgb(60, 64, 67); margin-bottom: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .TeNodb { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99 { background: rgb(255, 255, 255); display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: center; justify-content: center; cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AZW99 { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc { height: 64px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc .rNlsc { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc .O7pQ4 { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc .bRdBfe { width: 24px; height: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc .DcfYrb { width: 25px; height: 25px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.nhiZfc .kcuFCe { padding-left: 16px; padding-right: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd { height: 52px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd .rNlsc { font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; line-height: 1.25rem; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd .O7pQ4 { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; line-height: 1rem; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd .bRdBfe { width: 19px; height: 19px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd .DcfYrb { width: 20px; height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.XdSAtd .kcuFCe { padding-left: 12px; padding-right: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd { height: 44px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd .rNlsc { font-family: Roboto, Arial, sans-serif; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; line-height: 1.125; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd .O7pQ4 { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; line-height: 0.875rem; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd .bRdBfe { width: 17px; height: 17px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd .DcfYrb { width: 20px; height: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.HddOwd .kcuFCe { padding-left: 12px; padding-right: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.RDPZE { cursor: default; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.RDPZE .rNlsc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.RDPZE .G1zVib { color: rgb(60, 64, 67); opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AZW99.RDPZE .rNlsc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AZW99.RDPZE .G1zVib { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.RDPZE .p1rXue { opacity: 0.5; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.KKjvXb .s38Kwb { opacity: 1; transform: scale(1); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99:hover { background: rgba(10, 10, 10, 0.04); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AZW99:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.qs41qe { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .AZW99.qs41qe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .AZW99.FdSZEb { background-color: papayawhip; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .kcuFCe { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .r6EVzf { -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .uy8S0e { -webkit-box-flex: 1; flex: 1 1 auto; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .arWWkb { display: inline-flex; -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .CnoS1b { align-content: flex-start; -webkit-box-align: start; align-items: flex-start; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-flow: column nowrap; margin-left: 12px; margin-right: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pX5gAc { -webkit-box-flex: initial; flex: initial; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .rNlsc { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .PNwDub { color: rgb(60, 64, 67); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .PNwDub { color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .dUj0G { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-align: center; align-items: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .O7pQ4 { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .G1zVib { color: rgb(95, 99, 104); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .G1zVib { color: rgb(154, 160, 166); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .p1rXue { position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wRSMoe { height: inherit; width: inherit; position: relative; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .s38Kwb { background-color: rgb(26, 115, 232); border-radius: 50%; height: 100%; left: 0px; opacity: 0; outline: transparent solid 1px; position: absolute; top: 0px; transform: scale(0); transition: transform 0.15s ease-out 0s, -webkit-transform 0.15s ease-out 0s; width: 100%; display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .s38Kwb { background-color: rgb(138, 180, 248); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .GeKaSb { fill: rgb(255, 255, 255); display: inline-flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .GeKaSb { fill: rgb(32, 33, 36); }

@media (forced-colors: active) and (prefers-color-scheme: light) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .GeKaSb { filter: invert(1); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Hcawbb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; color: rgb(95, 99, 104); overflow: hidden; text-overflow: ellipsis; white-space: nowrap; display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .DcfYrb { margin-left: 16px; margin-right: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .DcfYrb[src=""] { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .S3hTZb { background-color: rgb(241, 243, 244); color: rgb(32, 33, 36); display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-align: center; align-items: center; margin-left: 8px; border-radius: 4px; outline: transparent solid 1px; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .S3hTZb.rNe0id { background-color: rgb(251, 188, 4); color: rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .nhiZfc .S3hTZb { height: 20px; min-width: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XdSAtd .S3hTZb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HddOwd .S3hTZb { height: 16px; min-width: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .nhiZfc .iHLOxc { width: 16px; height: 16px; margin-left: 2px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XdSAtd .iHLOxc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HddOwd .iHLOxc { width: 14px; height: 14px; margin-left: 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .R8dRld { max-width: 0px; overflow: hidden; transition: max-width 0.3s ease 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .S3hTZb:hover .R8dRld { max-width: 1000px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .xvZBXb { margin-left: 4px; margin-right: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .nhiZfc .xvZBXb { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0178571em; font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XdSAtd .xvZBXb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HddOwd .xvZBXb { font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.75rem; letter-spacing: 0.025em; font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .KMIgo { -webkit-box-align: center; align-items: center; display: flex; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .US5TTd { font-family: Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 400; color: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .US5TTd { color: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .l71Ouc { display: flex; -webkit-box-align: center; align-items: center; -webkit-box-pack: center; justify-content: center; background-color: rgb(241, 243, 244); border-radius: 50px; width: 32px; height: 32px; margin-left: 16px; margin-right: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .l71Ouc { background-color: rgba(241, 243, 244, 0.14); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .LYstE { fill: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .LYstE { fill: rgb(232, 234, 237); }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .LYstE { filter: brightness(0) invert(1); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc { background: none; border: none; border-radius: 50%; cursor: pointer; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc:hover { background-color: rgb(218, 220, 224); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .IYrrvc:hover { background-color: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc:active { background-color: rgb(189, 193, 198); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .IYrrvc:active { background-color: rgb(128, 134, 139); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.u3bW4e { background-color: rgb(218, 220, 224); outline: transparent solid 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .IYrrvc.u3bW4e { background-color: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.nhiZfc { height: 40px; padding: 8px; width: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.nhiZfc .ssmXx { height: 24px; width: 24px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.XdSAtd { height: 32px; padding: 6px; width: 32px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.XdSAtd .ssmXx { height: 20px; width: 20px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.HddOwd { height: 28px; padding: 5px; width: 28px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc.HddOwd .ssmXx { height: 18px; width: 18px; }

@media (forced-colors: active) and (prefers-color-scheme: dark) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IYrrvc .ssmXx { filter: brightness(0) invert(1); }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .L5nWEe { font-family: Roboto, Arial, sans-serif; font-size: 0.75rem; letter-spacing: 0.025em; background-color: rgb(60, 64, 67); color: rgb(241, 243, 244); border-radius: 5px; box-sizing: border-box; line-height: 16px; min-width: 40px; max-width: 200px; min-height: 24px; max-height: 40vh; overflow: hidden; padding: 4px 8px; position: fixed; outline: transparent solid 1px; text-align: center; font-weight: bold; width: max-content; z-index: 9; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .L5nWEe { background-color: rgb(60, 64, 67); color: rgb(232, 234, 237); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hxyQfd { -webkit-box-align: center; align-items: center; border-radius: 50%; cursor: pointer; display: flex; transition: transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hxyQfd:hover { background: rgba(10, 10, 10, 0.04); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .hxyQfd:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hxyQfd:active { background: rgba(10, 10, 10, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .hxyQfd:active { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hxyQfd.TICPrf { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .hxyQfd.TICPrf { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .hxyQfd.ReqAjb { transform: rotate(-180deg); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .e63afb { fill: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .e63afb { fill: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EhtNt { -webkit-box-align: center; align-items: center; border-radius: 50%; cursor: pointer; display: flex; transition: transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s, -webkit-transform 365ms cubic-bezier(0.4, 0, 0.2, 1) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EhtNt:hover { background: rgba(10, 10, 10, 0.04); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .EhtNt:hover { background: linear-gradient(0deg, rgba(232, 234, 237, 0.14), rgba(232, 234, 237, 0.14)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EhtNt:active { background: rgba(10, 10, 10, 0.12); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .EhtNt:active { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EhtNt.TICPrf { background: rgba(10, 10, 10, 0.12); outline: transparent solid 3px; outline-offset: -3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .EhtNt.TICPrf { background: linear-gradient(0deg, rgba(232, 234, 237, 0.19), rgba(232, 234, 237, 0.19)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .LGD9cb { fill: rgb(95, 99, 104); height: 16px; padding: 5px; width: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .LGD9cb { fill: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XhBoVe { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .XhBoVe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .a2oM9e { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-flow: row nowrap; padding-left: 16px; padding-right: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .TUsLr { color: rgb(95, 99, 104); font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.6875rem; letter-spacing: 0.0727273em; font-weight: 500; text-transform: uppercase; padding-bottom: 12px; padding-top: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .TUsLr { color: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .xvJ2yc { flex-shrink: initial; flex-basis: initial; -webkit-box-flex: 1; flex-grow: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .xAiMkd { -webkit-box-align: center; align-items: center; display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: normal; flex-direction: row; -webkit-box-pack: justify; justify-content: space-between; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .F2iRTc { -webkit-box-flex: initial; flex: initial; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .GZQpmf { -webkit-box-flex: initial; flex: initial; margin-left: 16px; margin-right: 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .RWYkoe { overflow: hidden; transform-origin: center top; transition: all 0.5s cubic-bezier(0.05, 0.7, 0.1, 1) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .RWYkoe.qAWA2 { height: 0px; transform: scaleY(0); transition: all 0.2s cubic-bezier(0.3, 0, 0.8, 0.15) 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .FDlMAe { background: rgb(255, 255, 255); color: rgb(95, 99, 104); font-family: Roboto, Arial, sans-serif; line-height: 1rem; font-size: 0.6875rem; letter-spacing: 0.0727273em; font-weight: 500; text-transform: uppercase; padding-bottom: 12px; padding-left: 16px; padding-top: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .FDlMAe { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); color: rgb(241, 243, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd { background: rgb(255, 255, 255); height: 100%; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; user-select: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .pIQtMd { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.JpY6Fd .L5WGxc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.JpY6Fd .zcyXfd { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.JpY6Fd .z7ZqLc { display: flex; -webkit-box-pack: center; justify-content: center; -webkit-box-align: center; align-items: center; height: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.JpY6Fd .z7ZqLc::before { -webkit-box-flex: 1; flex: 1 1 auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.JpY6Fd .z7ZqLc::after { -webkit-box-flex: 1; flex: 1 1 auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.Cn4kwe .L5WGxc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.Cn4kwe .z7ZqLc { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pIQtMd.Cn4kwe .zcyXfd { display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; -webkit-box-pack: start; justify-content: flex-start; -webkit-box-align: center; align-items: center; height: 100%; overflow: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .L5WGxc { height: 100%; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; overflow: hidden; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .z7ZqLc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .zcyXfd { display: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd { display: inline-block; height: 40px; position: relative; width: 40px; direction: ltr; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .FxUiNc { height: 0px; overflow: hidden; position: absolute; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .QPPI1e { width: 100%; height: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .QPPI1e { animation: 1568ms linear 0s infinite normal none running circular-progress-container-rotate; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .KLPWzf { height: 100%; opacity: 0; position: absolute; width: 100%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Y6U90b { border-color: rgb(66, 133, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .l36Xze { border-color: rgb(234, 67, 53); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .GybXwf { border-color: rgb(251, 188, 4); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .v5iurb { border-color: rgb(52, 168, 83); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .KLPWzf.Y6U90b { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-blue-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .KLPWzf.l36Xze { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-red-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .KLPWzf.GybXwf { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-yellow-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .KLPWzf.v5iurb { animation: 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-fill-unfill-rotate, 5332ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-green-fade-in-out; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .OEwgzc { position: absolute; box-sizing: border-box; top: 0px; left: 45%; width: 10%; height: 100%; overflow: hidden; border-color: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .OEwgzc .z58N3b { width: 1000%; left: -450%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tEVydc { display: inline-block; position: relative; width: 50%; height: 100%; overflow: hidden; border-color: inherit; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tEVydc .z58N3b { width: 200%; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .z58N3b { position: absolute; inset: 0px; box-sizing: border-box; height: 100%; border-width: 3px; border-style: solid; border-top-color: inherit; border-right-color: inherit; border-left-color: inherit; border-bottom-color: transparent; border-radius: 50%; animation: 0s ease 0s 1 normal none running none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tEVydc.A9Yu7d .z58N3b { border-right-color: transparent; transform: rotate(129deg); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tEVydc.scD29d .z58N3b { left: -100%; border-left-color: transparent; transform: rotate(-129deg); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .tEVydc.A9Yu7d .z58N3b { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-left-spin; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.qs41qe .tEVydc.scD29d .z58N3b { animation: 1333ms cubic-bezier(0.4, 0, 0.2, 1) 0s infinite normal both running circular-progress-right-spin; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .MFfTvd.sf4e6b .QPPI1e { animation: 1568ms linear 0s infinite normal none running circular-progress-container-rotate, 0.4s cubic-bezier(0.4, 0, 0.2, 1) 0s 1 normal none running circular-progress-fade-out; }

@-webkit-keyframes circular-progress-container-rotate { 
  100% { transform: rotate(1turn); }
}

@keyframes circular-progress-container-rotate { 
  100% { transform: rotate(1turn); }
}

@-webkit-keyframes circular-progress-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@keyframes circular-progress-fill-unfill-rotate { 
  12.5% { transform: rotate(135deg); }
  25% { transform: rotate(270deg); }
  37.5% { transform: rotate(405deg); }
  50% { transform: rotate(540deg); }
  62.5% { transform: rotate(675deg); }
  75% { transform: rotate(810deg); }
  87.5% { transform: rotate(945deg); }
  100% { transform: rotate(3turn); }
}

@-webkit-keyframes circular-progress-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@keyframes circular-progress-blue-fade-in-out { 
  0% { opacity: 0.99; }
  25% { opacity: 0.99; }
  26% { opacity: 0; }
  89% { opacity: 0; }
  90% { opacity: 0.99; }
  100% { opacity: 0.99; }
}

@-webkit-keyframes circular-progress-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@keyframes circular-progress-red-fade-in-out { 
  0% { opacity: 0; }
  15% { opacity: 0; }
  25% { opacity: 0.99; }
  50% { opacity: 0.99; }
  51% { opacity: 0; }
}

@-webkit-keyframes circular-progress-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@keyframes circular-progress-yellow-fade-in-out { 
  0% { opacity: 0; }
  40% { opacity: 0; }
  50% { opacity: 0.99; }
  75% { opacity: 0.99; }
  76% { opacity: 0; }
}

@-webkit-keyframes circular-progress-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes circular-progress-green-fade-in-out { 
  0% { opacity: 0; }
  65% { opacity: 0; }
  75% { opacity: 0.99; }
  90% { opacity: 0.99; }
  100% { opacity: 0; }
}

@-webkit-keyframes circular-progress-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@keyframes circular-progress-left-spin { 
  0% { transform: rotate(130deg); }
  50% { transform: rotate(-5deg); }
  100% { transform: rotate(130deg); }
}

@-webkit-keyframes circular-progress-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@keyframes circular-progress-right-spin { 
  0% { transform: rotate(-130deg); }
  50% { transform: rotate(5deg); }
  100% { transform: rotate(-130deg); }
}

@-webkit-keyframes circular-progress-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

@keyframes circular-progress-fade-out { 
  0% { opacity: 0.99; }
  100% { opacity: 0; }
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wZ7wOe { border: none; outline: none; overflow: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wZ7wOe::-webkit-scrollbar-thumb { background: rgb(221, 221, 221); border-width: 1px 4px; border-style: solid; border-color: white; border-radius: 8px; box-shadow: none; min-height: 40px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wZ7wOe::-webkit-scrollbar-thumb:active { background: rgb(95, 99, 104); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wZ7wOe:hover::-webkit-scrollbar-thumb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wZ7wOe::-webkit-scrollbar-thumb:hover { background: rgb(128, 134, 139); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HJOG0e { color: rgb(95, 99, 104); padding: 2em; text-align: center; -webkit-box-align: center; align-items: center; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .HJOG0e { color: rgb(154, 160, 166); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .E633ec { font-family: "Google Sans", Roboto, Arial, sans-serif; line-height: 1.5rem; font-size: 1rem; letter-spacing: 0.00625em; font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .LPP4B { font-family: Roboto, Arial, sans-serif; line-height: 1.25rem; font-size: 0.875rem; letter-spacing: 0.0142857em; font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .YlzPUb { color: inherit; text-decoration: underline; white-space: nowrap; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .OFaVze { border-width: 0px; box-shadow: rgba(60, 64, 67, 0.3) 0px 1px 3px 0px, rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; background: rgb(255, 255, 255); border-radius: 4px; display: flex; -webkit-box-orient: vertical; -webkit-box-direction: normal; flex-direction: column; outline: transparent solid 2px; overflow: hidden; padding-bottom: 8px; padding-top: 8px; position: absolute; user-select: none; z-index: 999999; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .OFaVze .VfPpkd-BFbNVe-bF1uUb { opacity: 0; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .aqWPhc .OFaVze { background: linear-gradient(0deg, rgba(232, 234, 237, 0.08), rgba(232, 234, 237, 0.08)), rgb(32, 33, 36); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-hFsbo-SmKAyb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-hFsbo-n0tgWb { display: none; }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-hFsbo-SmKAyb, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC-hFsbo-n0tgWb { height: 0px; position: absolute; width: 0px; }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb { border-top: none; border-bottom: 18px solid transparent; border-left: none; border-right: 18px solid rgb(255, 255, 255); left: -13px; top: 0px; }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-IIEkAe.wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb { border-right: 18px solid rgb(238, 238, 238); }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-n0tgWb { border-top: none; border-bottom: 24px solid transparent; border-left: none; border-right: 24px solid rgba(0, 0, 0, 0.133); left: -15px; top: -1px; z-index: -1; }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC > .wvGCSb-efwuC-hFsbo-SmKAyb, .wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-pnL5fc-auswjd.wvGCSb-efwuC > .wvGCSb-efwuC-hFsbo-n0tgWb { display: block; }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb.wvGCSb-JYA2rd-tSZMSb { border-right: 18px solid rgb(255, 255, 255); }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb.wvGCSb-JYA2rd-jf2N7b { border-right: 18px solid rgb(242, 242, 242); }

.wvGCSb-neVct-BvBYQ.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-efwuC .wvGCSb-efwuC-hFsbo-SmKAyb.wvGCSb-JYA2rd-dHwMxe { border-right: 18px solid rgb(66, 133, 244); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-Moncj-SmKAyb { border-top: 7px solid transparent; border-right: 8px solid rgb(255, 255, 255); border-bottom: 7px solid transparent; height: 0px; left: -6px; position: absolute; top: 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-YPqjbf-Moncj-n0tgWb { border-top: 7px solid transparent; border-right: 8px solid rgb(200, 200, 200); border-bottom: 7px solid transparent; height: 0px; left: -7px; position: absolute; top: 3px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .jCCvxc-hSRGPd-Sx9Kwc button.jCCvxc-hSRGPd-iib5kc-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .jCCvxc-hSRGPd-Sx9Kwc button.jCCvxc-hSRGPd-iib5kc-LgbsSe:hover { box-shadow: none; background-color: rgb(77, 144, 254); background-image: -webkit-gradient(linear, 0% 0%, 0% 100%, from(rgb(77, 144, 254)), to(rgb(71, 135, 237))); border: 1px solid rgb(48, 121, 237); color: rgb(255, 255, 255); }

.HB1eCd-HzV7m.VIpgJd-xl07Ob.VIpgJd-xl07Ob-RDtZlf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb, .HB1eCd-HzV7m.VIpgJd-xl07Ob.VIpgJd-xl07Ob-GP8zAc.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb { padding-left: 16px; }

.HB1eCd-HzV7m.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb { padding-left: 36px; }

.HB1eCd-HzV7m.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IyROMc-j7LFlb .VIpgJd-j7LFlb-MPu53c, .HB1eCd-HzV7m.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IyROMc-j7LFlb .VIpgJd-j7LFlb-Bz112c { left: 8px; }

.HB1eCd-HzV7m.VIpgJd-xl07Ob.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IyROMc-j7LFlb.VIpgJd-wQNmvb-gk6SMd { background-position: left 5px center; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.VIpgJd-xl07Ob .IyROMc-j7LFlb.VIpgJd-wQNmvb-gk6SMd { background-image: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m.VIpgJd-xl07Ob .IyROMc-j7LFlb.VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-MPu53c { background: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg") -62px -9766px no-repeat; height: 18px; width: 18px; top: 50%; margin-top: -9px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe { border: 1px solid transparent; border-radius: 4px; box-shadow: none; color: rgb(32, 33, 36); cursor: pointer; font-size: 14px; letter-spacing: 0.2px; padding: 4px 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-ZmdkE { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-FNFY6c { background-color: rgb(232, 240, 254); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe:hover:active { background-color: rgb(210, 227, 252); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-OWB6Me { color: rgb(154, 160, 166); background-color: white; cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .HB1eCd-xl07Ob-LgbsSe-FNFY6c-uFfGwd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .HB1eCd-xl07Ob-LgbsSe-FNFY6c-KLRBe { z-index: 1003; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe.HB1eCd-xl07Ob-LgbsSe-FNFY6c-uFfGwd { border-bottom-left-radius: 0px; border-bottom-right-radius: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob.HB1eCd-xl07Ob-M7EJ5d-LgbsSe-KLRBe { border-top-left-radius: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob.HB1eCd-xl07Ob-M7EJ5d-LgbsSe-uFfGwd { border-bottom-left-radius: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob { border: 1px solid transparent; border-radius: 4px; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; max-height: calc(100vh - 94px); overflow-y: auto; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob .VIpgJd-hEj1I-fFW7wc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob.HB1eCd-ex68ab { overflow: hidden; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob.HB1eCd-CtVXDf-YPIHXb-xl07Ob { overflow: visible; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ex68ab { max-height: unset; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-gqMrKb { border-top: 1px solid rgb(218, 220, 224); margin: 8px 0px 8px 36px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Y8b4pe .VIpgJd-gqMrKb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-vKt3Ub-zTETae-xl07Ob .VIpgJd-gqMrKb { margin-left: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-GP8zAc .VIpgJd-gqMrKb { margin-left: 13px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb { color: rgb(32, 33, 36); font-size: 14px; letter-spacing: 0.2px; line-height: 20px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob .VIpgJd-j7LFlb { padding: 6px 15px 6px 38px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob-GP8zAc .VIpgJd-j7LFlb { padding-left: 15px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob .IyROMc-j7LFlb .VIpgJd-j7LFlb-MPu53c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob .IyROMc-j7LFlb .VIpgJd-j7LFlb-Bz112c:not(.HB1eCd-QbdDtf-oKdM2c-Bz112c) { margin: 7px 8px 7px 12px; left: 0px; top: 0px; }

.HB1eCd-UMrnmb.HB1eCd-Guievd-WqyaDf.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-xl07Ob .IyROMc-j7LFlb .VIpgJd-j7LFlb-MPu53c { filter: invert(100%); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb .VIpgJd-j7LFlb-bN97Pc { min-height: 20px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb .VIpgJd-eKm5Fc-hFsbo { padding-top: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb .HB1eCd-INgbqf-WAutxc-OomVLb-xl07Ob-ij8cu, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb .HB1eCd-KVuj8d-Zr8acc-INgbqf-j7LFlb-ij8cu, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb .usbjsf-UmQjBf-F2hcT-nUpftc-xl07Ob-ibnC6b-ij8cu { color: rgb(95, 99, 104); font-size: 12px; line-height: 1; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q { border: none; background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-mZGCQb.VIpgJd-j7LFlb { padding-right: 10px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-ex68ab .VIpgJd-j7LFlb { padding-right: 48px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-bN97Pc { color: rgb(154, 160, 166) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-auswjd:hover:active { background-color: rgb(232, 234, 237); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-x29Bmf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-x29Bmf { color: rgb(128, 134, 139); font-weight: 500; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-CtVXDf-YPIHXb-xl07Ob-hFsbo-WgXLxe { border: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-QbdDtf-h0T7hb .VIpgJd-j7LFlb-Bz112c { top: auto; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-bN97Pc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-V67aGc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-x29Bmf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-sn54Q .VIpgJd-eKm5Fc-hFsbo, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-FNFY6c { forced-color-adjust: none; background-color: highlight !important; color: highlighttext !important; }
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe { border-color: canvas; }
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-loREFf .VIpgJd-bMcfAe-FNFY6c { border-color: highlight; }
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-bN97Pc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-V67aGc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-j7LFlb-x29Bmf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-OWB6Me .VIpgJd-eKm5Fc-hFsbo { color: graytext !important; }
}

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { opacity: 0.38; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar { height: 16px; overflow: visible; width: 16px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-button { height: 0px; width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track { background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 0px 0px 0px 4px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:horizontal { border-width: 4px 0px 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.1) 1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(0, 0, 0, 0.1) 0px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:active { background-color: rgba(0, 0, 0, 0.05); box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.2) 1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:horizontal:hover { box-shadow: rgba(255, 255, 255, 0.2) 0px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:active { background-color: rgba(255, 255, 255, 0.1); box-shadow: rgba(255, 255, 255, 0.25) 1px 0px 0px inset, rgba(255, 255, 255, 0.15) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:horizontal:active { box-shadow: rgba(255, 255, 255, 0.25) 0px 1px 0px inset, rgba(255, 255, 255, 0.15) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb { background-color: rgba(0, 0, 0, 0.2); background-clip: padding-box; border-style: solid; border-color: transparent; border-image: initial; border-width: 1px 1px 1px 6px; min-height: 28px; padding: 100px 0px 0px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb:horizontal { border-width: 6px 1px 1px; padding: 0px 0px 0px 100px; box-shadow: rgba(0, 0, 0, 0.1) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb:hover { background-color: rgba(0, 0, 0, 0.4); box-shadow: rgba(0, 0, 0, 0.25) 1px 1px 1px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb:active { background-color: rgba(0, 0, 0, 0.5); box-shadow: rgba(0, 0, 0, 0.35) 1px 1px 3px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb { background-color: rgba(255, 255, 255, 0.3); box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:horizontal { box-shadow: rgba(255, 255, 255, 0.15) 1px 1px 0px inset, rgba(255, 255, 255, 0.1) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:hover { background-color: rgba(255, 255, 255, 0.6); box-shadow: rgba(255, 255, 255, 0.37) 1px 1px 1px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-to915::-webkit-scrollbar-thumb:active { background-color: rgba(255, 255, 255, 0.75); box-shadow: rgba(255, 255, 255, 0.5) 1px 1px 3px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track { border-width: 0px 1px 0px 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track:horizontal { border-width: 6px 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-track:hover { background-color: rgba(0, 0, 0, 0.035); box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset, rgba(0, 0, 0, 0.07) -1px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G.tk3N6e-qrhCuc-to915::-webkit-scrollbar-track:hover { background-color: rgba(255, 255, 255, 0.07); box-shadow: rgba(255, 255, 255, 0.25) 1px 1px 0px inset, rgba(255, 255, 255, 0.15) -1px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-thumb { border-width: 0px 1px 0px 6px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-qrhCuc-xTH6G::-webkit-scrollbar-thumb:horizontal { border-width: 6px 0px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-corner { background: transparent; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body::-webkit-scrollbar-track-piece { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 0px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 0px 0px inset, rgba(0, 0, 0, 0.07) -1px 0px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body::-webkit-scrollbar-track-piece:horizontal { border-width: 3px 0px 0px; box-shadow: rgba(0, 0, 0, 0.14) 0px 1px 0px inset, rgba(0, 0, 0, 0.07) 0px -1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body::-webkit-scrollbar-thumb { border-width: 1px 1px 1px 5px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body::-webkit-scrollbar-thumb:horizontal { border-width: 5px 1px 1px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb body::-webkit-scrollbar-corner { background-clip: padding-box; background-color: rgb(245, 245, 245); border-style: solid; border-color: rgb(255, 255, 255); border-image: initial; border-width: 3px 0px 0px 3px; box-shadow: rgba(0, 0, 0, 0.14) 1px 1px 0px inset; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe-Kb3HCc { font-weight: normal; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-INgbqf-xl07Ob-LgbsSe { font-weight: 500; font-size: 12px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-editor, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-editor-container { background: rgb(248, 249, 250); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf #docs-editor, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf #docs-editor-container { background: rgb(249, 251, 253); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-MqDS2b-uoC0bf.HB1eCd-R1gDOc #docs-editor-container { background: rgb(255, 255, 255); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-AznF2e { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { font-weight: 400; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke { font-size: 22px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-F79BRe .VIpgJd-VgwJlc-PBWx0c, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-eLJrl { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-rugWtd-xGWjg, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-rugWtd-xGWjg:hover { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LR6Drb { font-weight: 500; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc { font-weight: 500; font-size: 12px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc { border-color: rgb(218, 220, 224) transparent; }

@media (forced-colors: active) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd.HB1eCd-EfADOe-VCkuzd { border: 1px solid canvastext; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd .tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border-color: canvastext canvas; }
  @supports (forced-color-adjust:none) {
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc-ez0xG, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe .tk3N6e-VCkuzd-jQ8oHc, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe .tk3N6e-VCkuzd-ez0xG { forced-color-adjust: none; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc { border-color: canvastext transparent; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG { border-color: canvas transparent; }
  .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-UMrnmb-EfADOe.tk3N6e-VCkuzd.tk3N6e-VCkuzd-EfADOe.HB1eCd-EfADOe-VCkuzd .tk3N6e-VCkuzd-hFsbo-hUbt4d.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG { border-color: canvastext transparent; }
}
}

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IyROMc-t6O8cf-r4nke-haAclf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .IyROMc-w3KqTd-r4nke-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-E90Ek-haAclf { font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-tCYPLb-LkdAo, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-tCYPLb-DbqQVb, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-jEqmyf-oPu43, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-k6D2ve-cXXICe-LYNcwc { background-color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-tCYPLb-i5vt6e, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-jEqmyf-VtOx3e, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-bwj4ec-VtOx3e { border-color: rgb(26, 115, 232); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-tCYPLb-DbqQVb { height: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); cursor: pointer; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-QDgCrf { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-NziyQe.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .usbjsf-OiiCO-PvRhvb-QKiGd.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-no16zc-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); cursor: pointer; border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-QDgCrf, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-QDgCrf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-QDgCrf { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HiaYvf-R5U1Nd-Of6OMd-S9gUrf-LgbsSe.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .pD2Zae-Irdsic-LgbsSe-haAclf .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-JEtDLd-ERydpb-haAclf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .h5F6zd-vWsuo .usbjsf-OiiCO-PvRhvb-htvI8d.VIpgJd-Kb3HCc-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; cursor: default; border: 1px solid rgb(241, 243, 244) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: white; color: rgb(26, 115, 232); border: 1px solid rgb(218, 220, 224) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:hover, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE { background: rgb(248, 251, 255); border: 1px solid rgb(204, 224, 252) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { background: rgb(233, 241, 254); border: 1px solid rgb(193, 216, 251) !important; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe { border: 1px solid highlight; }
}

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:hover:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { background: rgb(225, 236, 254); border: 1px solid rgb(187, 212, 251) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button:focus:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd { background: rgb(225, 236, 254); box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button[disabled], .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me { background: white; color: rgb(60, 64, 67); opacity: 0.38; border: 1px solid rgb(241, 243, 244) !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc { border-radius: 4px; box-shadow: none; box-sizing: border-box; font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-weight: 500; font-size: 14px; height: 36px; letter-spacing: 0.25px; line-height: 16px; padding: 9px 24px 11px; background: rgb(26, 115, 232); color: rgb(255, 255, 255); border: 1px solid transparent !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:hover, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE { color: rgb(255, 255, 255); background: rgb(43, 125, 233); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(80, 148, 237); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:hover:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE.tk3N6e-LgbsSe-XpnDCe { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 1px 3px 1px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc:focus:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-auswjd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-AHmuwe.tk3N6e-LgbsSe-auswjd { color: rgb(255, 255, 255); background: rgb(99, 160, 239); box-shadow: rgba(66, 133, 244, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc[disabled], .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { background: rgb(248, 249, 250); color: rgb(32, 33, 36); opacity: 0.62; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-n2to0e, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc { cursor: pointer; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-LgbsSe.VIpgJd-Kb3HCc-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc button[disabled], .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-ldDVFe-JIbuQc[disabled], .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me { cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .tk3N6e-y4JFTd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-y4JFTd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; color: rgb(60, 64, 67); padding: 1px 8px; font-size: 14px; height: 36px; margin: 8px 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc textarea.tk3N6e-y4JFTd { min-height: 36px; height: unset; padding: 7px 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc textarea.tk3N6e-y4JFTd { min-height: 52px; max-height: 52px; min-width: 100%; height: unset; padding: 7px 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-VCkuzd .tk3N6e-y4JFTd:focus { border: 2px solid rgb(26, 115, 232); box-shadow: none; padding: 0px 7px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc textarea.tk3N6e-y4JFTd:focus, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc textarea.tk3N6e-y4JFTd:focus { padding: 6px 7px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover { opacity: 1; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { background-color: transparent; border-radius: 50%; cursor: pointer; line-height: 18px; text-align: center; color: rgb(95, 99, 104); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: rgb(232, 234, 237); outline: none; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc { color: canvastext; }
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:hover, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: highlight; color: highlighttext; }
}

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-y4JFTd.EX2EHc-cwdWJf-rygyx { margin: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc.jcJzye-dZ8yzd-fFW7wc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF.tk3N6e-VCkuzd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Yygnk-uDEFge-V68bde.tk3N6e-VCkuzd { background: rgb(255, 255, 255); border: 1px solid transparent; border-radius: 8px; box-shadow: rgba(60, 64, 67, 0.15) 0px 4px 8px 3px; position: absolute; z-index: 1003; padding: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .fFW7wc.XKSfm-Sx9Kwc { padding: 0px; z-index: 1201; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc.jcJzye-dZ8yzd-fFW7wc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-bN97Pc, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-offline-optinpromo-description, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-offline-optinpromo-learn-more-container { color: rgb(60, 64, 67); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb #docs-offline-optinpromo-title { border-bottom: none; padding: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-r4nke-fmcmS { color: rgb(32, 33, 36); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 22px; font-weight: 400; line-height: 28px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd { display: flex; -webkit-box-orient: horizontal; -webkit-box-direction: reverse; flex-direction: row-reverse; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-McfNlf-c6xFrd { margin-top: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-PrY1nf-a3aHF-c6xFrd .tk3N6e-LgbsSe { cursor: pointer; margin-left: 16px; margin-right: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-NRdnKf-c6xFrd { display: flex; -webkit-box-pack: end; justify-content: flex-end; margin-top: 24px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button { margin: 0px 0px 0px 12px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd button:first-child { margin-left: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke { position: relative; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-fmcmS { display: inline-block; max-width: calc(100% - 32px); min-width: 200px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc { background-color: transparent; border-radius: 50%; cursor: pointer; height: 18px; line-height: 18px; padding: 7px; right: 0px; text-align: center; top: -3px; width: 18px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:hover { background-color: rgb(241, 243, 244); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:focus { background-color: rgb(232, 234, 237); outline: none; }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc:focus { border: 1px solid highlight; padding: 6px; }
}

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-Sx9Kwc .XKSfm-Sx9Kwc-r4nke-TvD9Pc::after { position: relative; right: 0px; top: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .HB1eCd-zPvuGf .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { height: 22px; width: 22px; border-radius: 50%; border: 1px solid rgb(218, 220, 224); margin: 0px; outline: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .HB1eCd-zPvuGf.VIpgJd-Kb3HCc-xl07Ob-LgbsSe { padding: 6px 0px 6px 6px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.VIpgJd-TUo6Hb-xJ5Hnf, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb div.XKSfm-Sx9Kwc-xJ5Hnf { background-color: rgb(0, 0, 0); left: 0px; position: absolute; top: 0px; z-index: 998; opacity: 0.6 !important; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track { box-shadow: none; margin: 0px 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-track:hover { box-shadow: none; background: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb { border-style: solid; border-color: transparent; border-width: 4px; background-color: rgb(218, 220, 224); border-radius: 8px; box-shadow: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb:hover { background-color: rgb(128, 134, 139); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb ::-webkit-scrollbar-thumb:active { background-color: rgb(95, 99, 104); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe { border: 1px solid rgb(218, 220, 224); border-radius: 4px; box-sizing: border-box; cursor: pointer; padding: 8px 6px 8px 8px; -webkit-box-align: center; align-items: center; background: none; color: rgb(60, 64, 67); display: inline-flex; -webkit-box-pack: justify; justify-content: space-between; outline: none; position: relative; width: unset; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { color: rgb(95, 99, 104); opacity: 0.38; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active { background-color: rgb(255, 255, 255); border: 1px solid transparent; box-shadow: rgba(60, 64, 67, 0.15) 0px 2px 6px 2px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE { background-color: rgba(60, 64, 67, 0.04); border: 1px solid rgb(218, 220, 224); box-shadow: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { background-color: rgba(60, 64, 67, 0.06); border: 1px solid rgb(218, 220, 224); }

@media screen and (forced-colors: active) {
  .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe { border: 1px solid highlight; }
}

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.04); border: 1px solid transparent; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-ZmdkE.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.06); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-XpnDCe.VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c { background-color: rgba(60, 64, 67, 0.08); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me { border: 1px solid rgb(218, 220, 224); box-shadow: none; cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { box-sizing: border-box; color: rgb(32, 33, 36); font-family: Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; height: 20px; line-height: 20px; max-width: 100%; overflow: hidden; text-overflow: ellipsis; white-space: nowrap; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-cHYyed { color: rgb(95, 99, 104); opacity: 0.38; cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { background: url("//ssl.gstatic.com/docs/common/material_common_sprite531_grey_medium.svg") -48px -12142px no-repeat; height: 18px; width: 18px; border: none; margin-top: 0px; position: relative; right: 0px; top: 0px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .HB1eCd-HzV7m-UMrnmb-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { opacity: 0.38; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-OWB6Me.VIpgJd-Kb3HCc-xl07Ob-LgbsSe:active { border: 1px solid rgb(218, 220, 224); cursor: default; box-shadow: none; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .Td0Hgc-PdaOHc-bMcfAe .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .EX2EHc-RbRzK-DpzZDb-bnBfGc-jXK9ad .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-FNFY6c .VIpgJd-Kb3HCc-xl07Ob-LgbsSe-j4gsHd { transform: rotate(180deg); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc .tk3N6e-Ru3Ixf-OWB6Me .tk3N6e-Ru3Ixf-V67aGc { color: rgb(95, 99, 104); opacity: 0.38; cursor: default; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-X3SwIb-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 14px; font-weight: 400; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-CJXtmf-Sx9Kwc .euCgFf-X3SwIb-haAclf { font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd { height: 40px; padding: 0px 16px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-X3SwIb-haAclf .tk3N6e-cXJiPb-TSZdd > span { display: flex; padding-top: 4px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-Bz112c { margin-right: 8px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-hSRGPd, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-hSRGPd:visited { color: rgb(26, 115, 232); font-family: "Google Sans", Roboto, RobotoDraft, Helvetica, Arial, sans-serif; font-size: 16px; margin-left: 80px; }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-hSRGPd:hover, .HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-hSRGPd:active { color: rgb(24, 90, 188); }

.HB1eCd-UMrnmb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .euCgFf-PLEiK-hSRGPd:disabled { color: rgb(26, 115, 232); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-LgbsSe { box-sizing: content-box; min-height: 0px; overflow: inherit; text-transform: none; transition: all 0s ease 0s; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c::before { border: 0px; border-radius: 0px; box-shadow: none; content: normal; height: auto; left: auto; margin: 0px; opacity: 1; position: static; top: auto; transition: all 0s ease 0s; width: auto; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c:hover::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c.tk3N6e-MPu53c-ZmdkE::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c:focus::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c.tk3N6e-MPu53c-XpnDCe::before { box-shadow: none; opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c:active::before, .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .tk3N6e-MPu53c.tk3N6e-MPu53c-auswjd::before { box-shadow: none; opacity: 1; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb { color: rgb(60, 64, 67); min-height: 0px; min-width: 0px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .VIpgJd-j7LFlb-bN97Pc { box-sizing: content-box; font-size: inherit; line-height: normal; min-height: 0px; padding: 0px; position: static; color: rgb(51, 51, 51); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.XKSfm-Sx9Kwc { border-radius: 0px; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb.XKSfm-Sx9Kwc { background: rgb(31, 31, 31); color: rgb(227, 227, 227); padding: 24px; border-radius: 8px; font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-size: 13px; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc { cursor: default; margin: 0px; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-TvD9Pc { display: none; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke { background-color: rgb(31, 31, 31); color: rgb(227, 227, 227); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 24px; line-height: 32px; margin: 0px 0px 24px; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-bN97Pc { background-color: rgb(31, 31, 31); }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { -webkit-box-pack: start; justify-content: flex-start; text-transform: none; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd { margin-top: 24px; display: flex; -webkit-box-pack: end; justify-content: flex-end; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button { min-height: 0px; text-transform: none; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button { margin: 0px 0px 0px 24px; line-height: 20px; border-radius: 100px; background: rgb(31, 31, 31); color: rgb(168, 199, 250); font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 500; font-size: 14px; border: none; transition: none 0s ease 0s; cursor: pointer; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button::before { border: none; box-shadow: none; transition: none 0s ease 0s; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button:hover { background: rgba(168, 199, 250, 0.08); color: rgb(168, 199, 250); border: none; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button:focus, .ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd > button:active { background: rgba(168, 199, 250, 0.12); color: rgb(168, 199, 250); border: none; outline: none; box-shadow: none; }

.wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS { color: inherit; font-size: inherit; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS { font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 24px; line-height: 32px; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled] { background: rgb(31, 31, 31); color: rgb(227, 227, 227); }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-tJHJj { font-family: "Google Sans", Roboto, Arial, sans-serif; font-style: normal; font-weight: 400; font-size: 16px; line-height: 24px; }

.ndfHFb-c4YZDc-uoC0bf .wvGCSb.wvGCSb.wvGCSb.wvGCSb.wvGCSb .wvGCSb-vhxNkb-h9d3hd { right: auto; color: rgb(168, 199, 250); }

sentinel { }
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/svg+xml
Content-Transfer-Encoding: binary
Content-Location: https://ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg

<?xml version="1.0" encoding="UTF-8"?>
<!DOCTYPE svg  PUBLIC '-//W3C//DTD SVG 1.1//EN'  'http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd'>
<svg width="31px" height="3834px" preserveAspectRatio="none" version="1.1" viewBox="0 0 31 3834" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
 <g transform="translate(0,1632)">
  <path d="M20 2H4c-1.1 0-2 .9-2 2v18l4-4h14c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 14H4V4h16v12zm-9-5H7V9h4V5h2v4h4v2h-4v4h-2v-4z"/>
 </g>
 <g transform="translate(0,2602)">
  <path d="M20 2H4c-1.1 0-2 .9-2 2v18l4-4h14c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 14H4V4h16v12zm-9-5H7V9h4V5h2v4h4v2h-4v4h-2v-4z" fill="#fff"/>
 </g>
 <g transform="translate(0,1816)" fill="#fff">
  <path d="m17.705 10.14-3.405-6.1401h-4.6l-6.1 11 2.1 4h8.1027c0.4644 0.8028 1.1094 1.488 1.8795 2h-9.9822c-0.7 0-1.4-0.4-1.8-1.1l-2.1-4c-0.3-0.6-0.3-1.3 0-1.9l6.2-11c0.3-0.6 1-1 1.7-1h4.6c0.7 0 1.4 0.4 1.8 1l3.9307 7.0882c-0.3348-0.058-0.6792-0.0882-1.0307-0.0882-0.4446 0-0.878 0.0484-1.295 0.1401z"/>
  <path d="m15.222 11.338-2.3225-3.9382h-1.8l-4.5 7.8 0.7 1.3h5.7205c-0.0136-0.1649-0.0205-0.3316-0.0205-0.5 0-0.5179 0.0656-1.0206 0.189-1.5h-3.889l2.7-4.8 1.83 3.2533c0.3651-0.6182 0.8378-1.1652 1.3925-1.6151z"/>
  <path d="m20 20v-3h3v-2h-3v-3h-2v3h-3v2h3v3h2z"/>
 </g>
 <g transform="translate(0,1448)" fill="#fff">
  <path d="m17.705 10.14-3.405-6.1401h-4.6l-6.1 11 2.1 4h8.1027c0.4644 0.8028 1.1094 1.488 1.8795 2h-9.9822c-0.7 0-1.4-0.4-1.8-1.1l-2.1-4c-0.3-0.6-0.3-1.3 0-1.9l6.2-11c0.3-0.6 1-1 1.7-1h4.6c0.7 0 1.4 0.4 1.8 1l3.9307 7.0882c-0.3348-0.058-0.6792-0.0882-1.0307-0.0882-0.4446 0-0.878 0.0484-1.295 0.1401z"/>
  <path d="m15.222 11.338-2.3225-3.9382h-1.8l-4.5 7.8 0.7 1.3h5.7205c-0.0136-0.1649-0.0205-0.3316-0.0205-0.5 0-0.5179 0.0656-1.0206 0.189-1.5h-3.889l2.7-4.8 1.83 3.2533c0.3651-0.6182 0.8378-1.1652 1.3925-1.6151z"/>
  <path d="m20 20v-3h3v-2h-3v-3h-2v3h-3v2h3v3h2z"/>
 </g>
 <g transform="translate(0,896)" fill="#fff">
  <path d="m17.705 10.14-3.405-6.1401h-4.6l-6.1 11 2.1 4h8.1027c0.4644 0.8028 1.1094 1.488 1.8795 2h-9.9822c-0.7 0-1.4-0.4-1.8-1.1l-2.1-4c-0.3-0.6-0.3-1.3 0-1.9l6.2-11c0.3-0.6 1-1 1.7-1h4.6c0.7 0 1.4 0.4 1.8 1l3.9307 7.0882c-0.3348-0.058-0.6792-0.0882-1.0307-0.0882-0.4446 0-0.878 0.0484-1.295 0.1401z"/>
  <path d="m15.222 11.338-2.3225-3.9382h-1.8l-4.5 7.8 0.7 1.3h5.7205c-0.0136-0.1649-0.0205-0.3316-0.0205-0.5 0-0.5179 0.0656-1.0206 0.189-1.5h-3.889l2.7-4.8 1.83 3.2533c0.3651-0.6182 0.8378-1.1652 1.3925-1.6151z"/>
  <path d="m20 20v-3h3v-2h-3v-3h-2v3h-3v2h3v3h2z"/>
 </g>
 <g transform="translate(0,2464)">
  <radialGradient id="svgid_1_" cx="-54.965" cy="277.45" r="72.073" gradientTransform="matrix(.09 .0525 -.052 .0909 25.385 -11.881)" gradientUnits="userSpaceOnUse">
   <stop stop-color="#0DA960" offset="0"/>
   <stop stop-color="#069B5A" offset="1"/>
  </radialGradient>
  <polygon points="4.175 21 0 13.693 8 0 12 7" fill="url(#svgid_1_)"/>
  <radialGradient id="svgid_2_" cx="45.038" cy="296.69" r="71.785" gradientTransform="matrix(.09 .0525 -.052 .0909 25.385 -11.881)" gradientUnits="userSpaceOnUse">
   <stop stop-color="#4387FD" offset="0"/>
   <stop stop-color="#3078F0" offset=".65"/>
   <stop stop-color="#2B72EA" offset=".9099"/>
   <stop stop-color="#286EE6" offset="1"/>
  </radialGradient>
  <polygon points="4.175 21 8 14 24 14 19.825 21" fill="url(#svgid_2_)"/>
  <radialGradient id="svgid_3_" cx="11.704" cy="200.89" r="81.652" gradientTransform="matrix(.09 .0525 -.052 .0909 25.385 -11.881)" gradientUnits="userSpaceOnUse">
   <stop stop-color="#FFD24D" offset="0"/>
   <stop stop-color="#F6C338" offset="1"/>
  </radialGradient>
  <polygon points="24 14 16 14 8 0 16 0" fill="url(#svgid_3_)"/>
  <polygon points="12 14 8 14 10 11 4.175 21" fill="#231F20" opacity=".08"/>
  <polygon points="16 14 24 14 14 10" fill="#231F20" opacity=".08"/>
  <polygon points="10.175 10.5 12 7.307 7.824 0" fill="#231F20" opacity=".08"/>
  <radialGradient id="svgid_4_" cx="16.564" cy="7.6699" r="108.01" gradientTransform="matrix(.1039 0 0 .105 10.279 9.6947)" gradientUnits="userSpaceOnUse">
   <stop stop-color="#fff" stop-opacity=".1" offset="0"/>
   <stop stop-color="#fff" stop-opacity=".091" offset=".0896"/>
   <stop stop-color="#fff" stop-opacity="0" offset="1"/>
  </radialGradient>
  <path d="M24,13.693L16.175,0H7.824L0,13.693L4.175,21l15.65,0L24,13.693L24,13.693z M12,7.307l3.65,6.387 h-7.3L12,7.307z" fill="url(#svgid_4_)"/>
 </g>
 <g transform="translate(0,816)">
  <g fill="#fff">
   <path d="M8.214,16.2H6.5c-0.939,0-1.7-0.762-1.7-1.7s0.761-1.7,1.7-1.7h1.714c0.364,0,0.593,0.173,0.786,0.45h1     C9.707,12.541,8.947,12,8.214,12H6.5C5.118,12,4,13.12,4,14.5S5.118,17,6.5,17h1.714c0.733,0,1.493-0.541,1.786-1.25H9     C8.807,16.027,8.578,16.2,8.214,16.2z"/>
   <path d="M7,14.499C7,14.775,7.225,15,7.5,15h6c0.275,0,0.5-0.225,0.5-0.501S13.775,14,13.5,14h-6     C7.225,14,7,14.223,7,14.499z"/>
   <path d="m14.5 12h-1.715c-0.732 0-1.492 0.541-1.785 1.25h1c0.193-0.277 0.422-0.45 0.785-0.45h1.715c0.939 0 1.7 0.762 1.7 1.7s-0.761 1.7-1.7 1.7h-1.715c-0.363 0-0.592-0.173-0.785-0.45h-1c0.293 0.709 1.053 1.25 1.785 1.25h1.715c1.382 0 2.49-1.12 2.49-2.5s-1.108-2.5-2.49-2.5z"/>
   <path d="m11 7v-4h-5v8h9v-4h-4zm-3 2h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm2 4h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm2 4h-1v-1h1v1zm2 0h-1v-1h1v1z"/>
  </g>
 </g>
 <g transform="translate(0,736)">
  <g fill="#fff">
   <path d="m8.214 16.2h-1.714c-0.939 0-1.7-0.762-1.7-1.7s0.761-1.7 1.7-1.7h1.714c0.364 0 0.593 0.173 0.786 0.45h1c-0.293-0.709-1.053-1.25-1.786-1.25h-1.714c-1.382 0-2.5 1.12-2.5 2.5s1.118 2.5 2.5 2.5h1.714c0.733 0 1.493-0.541 1.786-1.25h-1c-0.193 0.277-0.422 0.45-0.786 0.45z"/>
   <path d="m7 14.499c0 0.276 0.225 0.501 0.5 0.501h6c0.275 0 0.5-0.225 0.5-0.501s-0.225-0.499-0.5-0.499h-6c-0.275 0-0.5 0.222-0.5 0.499z"/>
   <path d="m14.5 12h-1.715c-0.732 0-1.492 0.541-1.785 1.25h1c0.193-0.277 0.422-0.45 0.785-0.45h1.715c0.939 0 1.7 0.762 1.7 1.7s-0.761 1.7-1.7 1.7h-1.715c-0.363 0-0.592-0.173-0.785-0.45h-1c0.293 0.709 1.053 1.25 1.785 1.25h1.715c1.382 0 2.49-1.12 2.49-2.5s-1.108-2.5-2.49-2.5z"/>
   <path d="m11 7v-2h-5v6h9v-4h-4zm-3 2h-1v-1h1v1zm0-2h-1v-1h1v1zm2 2h-1v-1h1v1zm0-2h-1v-1h1v1zm2 2h-1v-1h1v1zm2 0h-1v-1h1v1z"/>
  </g>
 </g>
 <g transform="translate(0,3634)">
  <path d="m4 16v6h16v-6c0-1.1-0.9-2-2-2h-12c-1.1 0-2 0.9-2 2zm14 2h-12v-2h12v2zm-6-16c-2.76 0-5 2.24-5 5l5 7 5-7c0-2.76-2.24-5-5-5zm0 9-3-4c0-1.66 1.34-3 3-3s3 1.34 3 3l-3 4z"/>
 </g>
 <g transform="translate(0,2544)">
  <path d="m4 16v6h16v-6c0-1.1-0.9-2-2-2h-12c-1.1 0-2 0.9-2 2zm14 2h-12v-2h12v2zm-6-16c-2.76 0-5 2.24-5 5l5 7 5-7c0-2.76-2.24-5-5-5zm0 9-3-4c0-1.66 1.34-3 3-3s3 1.34 3 3l-3 4z" fill="#174ea6"/>
 </g>
 <g transform="translate(0,2850)">
  <path d="m4 16v6h16v-6c0-1.1-0.9-2-2-2h-12c-1.1 0-2 0.9-2 2zm14 2h-12v-2h12v2zm-6-16c-2.76 0-5 2.24-5 5l5 7 5-7c0-2.76-2.24-5-5-5zm0 9-3-4c0-1.66 1.34-3 3-3s3 1.34 3 3l-3 4z" fill="#fff"/>
 </g>
 <g transform="translate(0,936)" stroke="#FFF">
  <polygon points="5 12 8 12 14 6 14 22 8 16 5 16" fill="#FFF" stroke-linejoin="round" stroke-width="2.2"/>
  <path d="m17.5 11c1.5 1 1.5 4.5 0 5.5" fill="none" stroke-linecap="round" stroke-width="1.5"/>
  <path d="m19 9c3 1.5 3 8.5 0 10" fill="none" stroke-linecap="round" stroke-width="1.5"/>
  <path d="m21 7c4 2 4 12 0 14" fill="none" stroke-linecap="round" stroke-width="1.5"/>
 </g>
 <g transform="translate(0,3794)" stroke="#FFF">
  <polygon points="5 12 8 12 14 6 14 22 8 16 5 16" fill="#FFF" stroke-linejoin="round" stroke-width="2.2"/>
  <path d="m17.5 11c1.5 1 1.5 4.5 0 5.5" fill="none" stroke-linecap="round" stroke-width="1.5"/>
 </g>
 <g transform="translate(0,2810)" stroke="#FFF">
  <polygon points="5 12 8 12 14 6 14 22 8 16 5 16" fill="#FFF" stroke-linejoin="round" stroke-width="2.2"/>
  <path d="m17.5 11c1.5 1 1.5 4.5 0 5.5" fill="none" stroke-linecap="round" stroke-width="1.5"/>
  <path d="m19 9c3 1.5 3 8.5 0 10" fill="none" stroke-linecap="round" stroke-width="1.5"/>
 </g>
 <g transform="translate(0,1408)" fill="#fff">
  <path d="M5,17.1h1.134L15.1,8.134V6c0-0.445-0.268-0.846-0.679-1.016c-0.411-0.172-0.884-0.077-1.199,0.238 L7.544,10.9H5c-0.607,0-1.1,0.493-1.1,1.1v4C3.9,16.607,4.393,17.1,5,17.1z"/>
  <path d="M10.004,19.559l3.218,3.219C13.433,22.988,13.714,23.1,14,23.1c0.142,0,0.285-0.027,0.421-0.083 C14.832,22.846,15.1,22.445,15.1,22v-7.537L10.004,19.559z"/>
  <path d="m5.088 22.354 14.314-14.313c8e-3 -7e-3 0.018-0.01 0.025-0.017 0.271-0.295 0.267-0.75-0.019-1.035-0.289-0.293-0.759-0.292-1.052-5e-3 -0.012 0.014-0.017 0.031-0.029 0.044l-14.314 14.313c-2e-3 2e-3 -5e-3 3e-3 -7e-3 5e-3 -0.255 0.295-0.252 0.736 0.027 1.016 0.287 0.286 0.745 0.288 1.04 0.016 6e-3 -8e-3 8e-3 -0.018 0.015-0.024z"/>
 </g>
 <g transform="translate(0,2344)" fill="#FFF" stroke="#FFF" stroke-linejoin="round" stroke-width="3">
  <rect x="6" y="7" width="3" height="14"/>
  <rect x="14" y="7" width="3" height="14"/>
 </g>
 <g transform="translate(0,3386)">
  <polygon points="6 7 6 21 17 14" fill="#FFF" stroke="#FFF" stroke-linejoin="round" stroke-width="3"/>
 </g>
 <g transform="translate(0,1080)">
  <polygon points="12.723 15 8 11.048 12.713 7 14 8.408 10.947 11.029 13.99 13.576"/>
 </g>
 <g transform="translate(0,1240)">
  <path d="m12 2-11 19h22l-11-19zm0 16c-0.55 0-1-0.45-1-1s0.45-1 1-1 1 0.45 1 1-0.45 1-1 1zm-1-3v-5h2v5h-2z" enable-background="new"/>
 </g>
 <g transform="translate(0,88)">
  <path d="M22 9.24l-7.19-.62L12 2 9.19 8.63 2 9.24l5.46 4.73L5.82 21 12 17.27 18.18 21l-1.63-7.03L22 9.24zM12 15.4l-3.76 2.27 1-4.28-3.32-2.88 4.38-.38L12 6.1l1.71 4.04 4.38.38-3.32 2.88 1 4.28L12 15.4z"/>
 </g>
 <g transform="translate(0,1488)">
  <path d="M22 9.24l-7.19-.62L12 2 9.19 8.63 2 9.24l5.46 4.73L5.82 21 12 17.27 18.18 21l-1.63-7.03L22 9.24zM12 15.4l-3.76 2.27 1-4.28-3.32-2.88 4.38-.38L12 6.1l1.71 4.04 4.38.38-3.32 2.88 1 4.28L12 15.4z" fill="#fff"/>
 </g>
 <g transform="translate(0)">
  <g fill="#fff">
   <path d="m8.67 17.76h-1.645c-0.432-3.122-2.899-5.592-6.025-6.027v-1.633c4.024 0.449 7.217 3.638 7.67 7.66zm-2.86 0h-1.651c-0.371-1.559-1.596-2.786-3.159-3.155v-1.64c2.456 0.412 4.393 2.345 4.81 4.795zm-2.922 0h-1.888v-1.884c0.886 0.305 1.582 1.002 1.888 1.884z"/>
   <path d="M10.082,16.651c-0.106-0.508-0.252-1.006-0.431-1.49h8.856V4.729l-14.9-0.005v4.395     C3.128,8.94,2.628,8.795,2.118,8.691V3.24H20v13.411H10.082z"/>
  </g>
 </g>
 <g transform="translate(0,1976)">
  <g>
   <path d="m8.67 17.76h-1.645c-0.432-3.122-2.899-5.592-6.025-6.027v-1.633c4.024 0.449 7.217 3.638 7.67 7.66zm-2.86 0h-1.651c-0.371-1.559-1.596-2.786-3.159-3.155v-1.64c2.456 0.412 4.393 2.345 4.81 4.795zm-2.922 0h-1.888v-1.884c0.886 0.305 1.582 1.002 1.888 1.884z"/>
   <path d="M10.082,16.651c-0.106-0.508-0.252-1.006-0.431-1.49h8.856V4.729l-14.9-0.005v4.395     C3.128,8.94,2.628,8.795,2.118,8.691V3.24H20v13.411H10.082z"/>
  </g>
 </g>
 <g transform="translate(0,1528)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M20 11H7.83l5.59-5.59L12 4l-8 8 8 8 1.41-1.41L7.83 13H20v-2z" fill="#fff"/>
 </g>
 <g transform="translate(0,3178)">
  <path d="M19 6.41L17.59 5 12 10.59 6.41 5 5 6.41 10.59 12 5 17.59 6.41 19 12 13.41 17.59 19 19 17.59 13.41 12z" fill="#fff"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1160)">
  <path d="M19 6.41L17.59 5 12 10.59 6.41 5 5 6.41 10.59 12 5 17.59 6.41 19 12 13.41 17.59 19 19 17.59 13.41 12z" fill="#174ea6"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1120)">
  <path d="M19 6.41L17.59 5 12 10.59 6.41 5 5 6.41 10.59 12 5 17.59 6.41 19 12 13.41 17.59 19 19 17.59 13.41 12z" fill="#5f6368"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,3570)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M19 6.41L17.59 5 12 10.59 6.41 5 5 6.41 10.59 12 5 17.59 6.41 19 12 13.41 17.59 19 19 17.59 13.41 12 19 6.41z"/>
 </g>
 <g transform="translate(0,2642)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M21.99 4c0-1.1-.89-2-1.99-2H4c-1.1 0-2 .9-2 2v12c0 1.1.9 2 2 2h14l4 4-.01-18zM17 11h-4v4h-2v-4H7V9h4V5h2v4h4v2z"/>
 </g>
 <g transform="translate(0,40)" fill="#5F6368">
  <path d="m6.8285 4-2-2h15.172c1.1 0 1.99 0.9 1.99 2l0.0095 15.171-3.171-3.171h1.1715v-12h-13.172z"/>
  <path d="m8.8285 6h9.1715v2h-7.1715l-2-2z"/>
  <path d="m11.828 9h6.1715v2h-4.1715l-2-2z"/>
  <path d="m14.828 12h3.1715v2h-1.1715l-2-2z"/>
  <path d="m2.1005 2.1005-1.4142 1.4142 1.3137 1.3137v11.172c0 1.1 0.9 2 2 2h11.172l5.3137 5.3137 1.4142-1.4142-19.799-19.799zm1.8995 13.9v-9.1716l2.1716 2.1716h-0.17164v2h2.1716l1 1h-3.1716v2h5.1716l2 2h-9.1716z" clip-rule="evenodd" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,1304)">
  <mask id="mask2" x="4" y="2" width="16" height="20" mask-type="alpha" maskUnits="userSpaceOnUse">
   <path d="m12 2 8 3.64v5.45c0 5.05-3.4132 9.76-8 10.91-4.5868-1.15-8-5.86-8-10.91v-5.45l8-3.64zm0 2.1891-6.044 2.75v4.1509c0 3.9892 2.5975 7.7144 6.044 8.8336 3.4465-1.1192 6.044-4.8444 6.044-8.8336v-4.1509l-6.044-2.75zm0 3.8109c1.1046 0 2 0.87056 2 1.9444 0 0.73016-0.414 1.3664-1.0262 1.6988l0.6902 3.3568h-3.2l0.6796-3.2979c-0.6761-0.3119-1.1436-0.9817-1.1436-1.7577 0-1.0739 0.8954-1.9444 2-1.9444z" fill="#fff"/>
  </mask>
  <g mask="url(#mask2)">
   <rect width="24" height="24" fill="#5F6368"/>
  </g>
 </g>
 <g transform="translate(0,3338)">
  <mask id="mask1" x="4" y="2" width="16" height="20" mask-type="alpha" maskUnits="userSpaceOnUse">
   <path d="m12 2 8 3.64v5.45c0 5.05-3.4132 9.76-8 10.91-4.5868-1.15-8-5.86-8-10.91v-5.45l8-3.64zm0 2.1891-6.044 2.75v4.1509c0 3.9892 2.5975 7.7144 6.044 8.8336 3.4465-1.1192 6.044-4.8444 6.044-8.8336v-4.1509l-6.044-2.75zm0 3.8109c1.1046 0 2 0.87056 2 1.9444 0 0.73016-0.414 1.3664-1.0262 1.6988l0.6902 3.3568h-3.2l0.6796-3.2979c-0.6761-0.3119-1.1436-0.9817-1.1436-1.7577 0-1.0739 0.8954-1.9444 2-1.9444z" fill="#fff"/>
  </mask>
  <g mask="url(#mask1)">
   <path d="M24 0H0V24H24V0Z" fill="#fff"/>
  </g>
 </g>
 <g transform="translate(0,2584)">
  <path d="m11.25 2.25v0.75h3.75v1.5h-0.75v9.75c0 0.825-0.675 1.5-1.5 1.5h-7.5c-0.825 0-1.5-0.675-1.5-1.5v-9.75h-0.75v-1.5h3.75v-0.75h4.5zm-6 12h7.5v-9.75h-7.5v9.75zm1.5-8.25h1.5v6.75h-1.5v-6.75zm4.5 0h-1.5v6.75h1.5v-6.75z" clip-rule="evenodd" fill="#fff" fill-rule="evenodd"/>
  <mask id="mask0" x="3" y="2" width="12" height="14" mask-type="alpha" maskUnits="userSpaceOnUse">
   <path d="m11.25 2.25v0.75h3.75v1.5h-0.75v9.75c0 0.825-0.675 1.5-1.5 1.5h-7.5c-0.825 0-1.5-0.675-1.5-1.5v-9.75h-0.75v-1.5h3.75v-0.75h4.5zm-6 12h7.5v-9.75h-7.5v9.75zm1.5-8.25h1.5v6.75h-1.5v-6.75zm4.5 0h-1.5v6.75h1.5v-6.75z" clip-rule="evenodd" fill="#fff" fill-rule="evenodd"/>
  </mask>
  <g mask="url(#mask0)">
   <path d="M0 0H18V18H0V0Z" clip-rule="evenodd" fill="#fff" fill-rule="evenodd"/>
  </g>
 </g>
 <g transform="translate(0,2890)">
  <path d="M6 19c0 1.1.9 2 2 2h8c1.1 0 2-.9 2-2V7H6v12zM19 4h-3.5l-1-1h-5l-1 1H5v2h14V4z"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1712)">
  <path d="M11 17h2v-6h-2v6zm1-15C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zM11 9h2V7h-2v2z"/>
 </g>
 <g transform="translate(0,208)">
  <path d="M11 17h2v-6h-2v6zm1-15C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zM11 9h2V7h-2v2z" fill="#fff"/>
 </g>
 <g transform="translate(0,1264)">
  <path d="m11 9v-4h-7v11h13v-7h-6zm-4 5h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm2 6h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm0-2h-1v-1h1v1zm4 6h-1v-1h1v1zm0-2h-1v-1h1v1zm2 2h-1v-1h1v1zm0-2h-1v-1h1v1z" fill="#fff"/>
 </g>
 <g transform="translate(0,2384)">
  <path d="M4 15h2v3h12v-3h2v3c0 1.1-.9 2-2 2H6c-1.1 0-2-.9-2-2m11.59-8.41L13 12.17V4h-2v8.17L8.41 9.59 7 11l5 5 5-5-1.41-1.41z" fill="#fff"/>
 </g>
 <g transform="translate(0,632)">
  <path d="M4 15h2v3h12v-3h2v3c0 1.1-.9 2-2 2H6c-1.1 0-2-.9-2-2m11.59-8.41L13 12.17V4h-2v8.17L8.41 9.59 7 11l5 5 5-5-1.41-1.41z"/>
 </g>
 <g transform="translate(0,328)">
  <path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm-8.5 11l-1.1-2.14 2.84-4.96 1.5 2.66L12.25 17h-.75zm6.8 0h-5.55l1.4-2.5h5.11l.26.46L18.3 17zm-4.55-8h2.39l2.84 5h-2.93l-2.56-4.54.26-.46z" fill="#fff"/>
 </g>
 <g transform="translate(0,672)">
  <path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm-8.5 11l-1.1-2.14 2.84-4.96 1.5 2.66L12.25 17h-.75zm6.8 0h-5.55l1.4-2.5h5.11l.26.46L18.3 17zm-4.55-8h2.39l2.84 5h-2.93l-2.56-4.54.26-.46z"/>
 </g>
 <g transform="translate(0,288)">
  <path d="M3 17.25V21h3.75L17.81 9.94l-3.75-3.75L3 17.25zM20.71 7.04c.39-.39.39-1.02 0-1.41l-2.34-2.34c-.39-.39-1.02-.39-1.41 0l-1.83 1.83 3.75 3.75 1.83-1.83z" fill="#fff"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,3466)">
  <polygon points="21 10 31 10 21 0" fill="#bbb"/>
  <defs>
   <filter id="Adobe_OpacityMaskFilter" x="21" y="0" width="10" height="10" filterUnits="userSpaceOnUse">
    <feColorMatrix color-interpolation-filters="sRGB" result="source" values="-1 0 0 0 1  0 -1 0 0 1  0 0 -1 0 1  0 0 0 1 0"/>
   </filter>
  </defs>
  <mask id="SVGID_1_" x="21" y="0" width="10" height="10" maskUnits="userSpaceOnUse">
   <g filter="url(#Adobe_OpacityMaskFilter)">
    <image transform="translate(19 -1.9995)" width="14" height="14" overflow="visible" xlink:href="data:image/jpeg;base64,/9j/4AAQSkZJRgABAgEASABIAAD/7AARRHVja3kAAQAEAAAAHgAA/+4AIUFkb2JlAGTAAAAAAQMAEAMCAwYAAAGAAAABlwAAAeb/2wCEABALCwsMCxAMDBAXDw0PFxsUEBAUGx8XFxcXFx8eFxoaGhoXHh4jJSclIx4vLzMzLy9AQEBAQEBAQEBAQEBAQEABEQ8PERMRFRISFRQRFBEUGhQWFhQaJhoaHBoa JjAjHh4eHiMwKy4nJycuKzU1MDA1NUBAP0BAQEBAQEBAQEBAQP/CABEIAA4ADgMBIgACEQEDEQH/ xABzAAEBAAAAAAAAAAAAAAAAAAAGBQEBAAAAAAAAAAAAAAAAAAAAABAAAgMBAAAAAAAAAAAAAAAAAAQBBQYDEQACAQEGBwEAAAAAAAAAAAABAgMEABESIhMFECExQaEyciMSAQAAAAAAAAAAAAAAAAAA AAD/2gAMAwEAAhEDEQAAADEZ2aP/2gAIAQIAAQUAP//aAAgBAwABBQA//9oACAEBAAEFAOWadZpDJvabhSyxM33/2gAIAQICBj8Af//aAAgBAwIGPwB//9oACAEBAQY/ABu9KpkVSwljHNrlJF68Am37alXR4n/Vpo4+5xZXYGyzCkjEokzU2oumZPv16+bf/9k="></image>
   </g>
  </mask>
  <g mask="url(#SVGID_1_)" opacity=".17">
   <polygon points="21 10 31 10 21 0"/>
  </g>
  <path d="M20,11V0H3C1.344,0,0,1.344,0,3v31c0,1.657,1.344,3,3,3h25c1.657,0,3-1.343,3-3V11H20z M9,12     c1.657,0,3,1.343,3,3s-1.343,3-3,3s-3-1.343-3-3S7.344,12,9,12z M22.153,30c-1.383-2.048-3.96-3.429-6.919-3.429     S9.698,27.953,8.315,30C7.209,30,7,29.143,6,28.287C8,25.714,10.572,23,15.234,23S22,25.714,24,28.287     C23,29.143,23.361,30,22.153,30z M21,18c-1.656,0-3-1.343-3-3s1.344-3,3-3s3,1.343,3,3S22.657,18,21,18z" fill="#C9C9C9"/>
  <defs>
   <filter id="Adobe_OpacityMaskFilter_1_" x="0" y="0" width="31" height="37" filterUnits="userSpaceOnUse">
    <feColorMatrix color-interpolation-filters="sRGB" result="source" values="-1 0 0 0 1  0 -1 0 0 1  0 0 -1 0 1  0 0 0 1 0"/>
   </filter>
  </defs>
  <mask id="SVGID_2_" x="0" y="0" width="31" height="37" maskUnits="userSpaceOnUse">
   <g filter="url(#Adobe_OpacityMaskFilter_1_)">
    <image transform="translate(-1.9995 -1.9995)" width="35" height="41" overflow="visible" xlink:href="data:image/jpeg;base64,/9j/4AAQSkZJRgABAgEASABIAAD/7AARRHVja3kAAQAEAAAAHgAA/+4AIUFkb2JlAGTAAAAAAQMAEAMCAwYAAAG6AAACIAAAAuj/2wCEABALCwsMCxAMDBAXDw0PFxsUEBAUGx8XFxcXFx8eFxoaGhoXHh4jJSclIx4vLzMzLy9AQEBAQEBAQEBAQEBAQEABEQ8PERMRFRISFRQRFBEUGhQWFhQaJhoaHBoa JjAjHh4eHiMwKy4nJycuKzU1MDA1NUBAP0BAQEBAQEBAQEBAQP/CABEIACkAIwMBIgACEQEDEQH/ xACMAAACAwEBAAAAAAAAAAAAAAAABgIEBwUDAQEAAAAAAAAAAAAAAAAAAAAAEAABBAEDBAMAAAAAAAAAAAAFAgMEBgEAFAcQIDATERIXEQACAQMCAwMNAQAAAAAAAAABAhEAMQMhElETBLEihBAgQWFx gaEyQoKSFEQFEgEAAAAAAAAAAAAAAAAAAAAw/9oADAMBAAIRAxEAAADksPmyGeK+koZSJhoHQpVBjgtORlJIOw0ZWGs0c0C4Uw//2gAIAQIAAQUA8P8A/9oACAEDAAEFAPD/AP/aAAgBAQABBQCsVaOZY/Nx/wAWirshmenHjyGh0OyCpsvkdaMw2xM11r1L1QY24GC6YyMLWWuMH0prrI4R9Ma49e9Q0nPsRkhtbeKViauYD1Uz8QZHZuYJvK7yDVgjcxbsXco7v//aAAgBAgIGPwAf/9oACAEDAgY/AB//2gAIAQEBBj8A5uQm5BgkWr5m/I0MmMm4Gpm/ldnMAM3bR6PBmVswmVBE6aGkxlgrFhEmJjWucigpEzNW +rZ91OkwCWHxpv8AQOcmSxCmI7xnhWJRm2NjM92OEemjhB3nGsbjc6V4zbTm8Fu2nwdAH6fBiYqXII3EcJFqHVc09Sq6tjOkiv2MiFGdJKsCDbga8dRx53CySYPrNbt6Am9qg5FPtNNhw5F1EAA1f+jm+7zv/9k="></image>
   </g>
  </mask>
  <g mask="url(#SVGID_2_)" opacity=".15">
   <path d="M20,11V0H3C1.344,0,0,1.344,0,3v31c0,1.657,1.344,3,3,3h25c1.657,0,3-1.343,3-3V11H20z M9,12c1.657,0,3,1.343,3,3     s-1.343,3-3,3s-3-1.343-3-3S7.344,12,9,12z M22.153,30c-1.383-2.048-3.96-3.429-6.919-3.429S9.698,27.953,8.315,30     C7.209,30,7,29.143,6,28.287C8,25.714,10.572,23,15.234,23S22,25.714,24,28.287C23,29.143,23.361,30,22.153,30z M21,18     c-1.656,0-3-1.343-3-3s1.344-3,3-3s3,1.343,3,3S22.657,18,21,18z"/>
  </g>
 </g>
 <g transform="translate(0,2240)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M11 15h2v2h-2v-2zm0-8h2v6h-2V7zm.99-5C6.47 2 2 6.48 2 12s4.47 10 9.99 10C17.52 22 22 17.52 22 12S17.52 2 11.99 2zM12 20c-4.42 0-8-3.58-8-8s3.58-8 8-8 8 3.58 8 8-3.58 8-8 8z" fill="#D93025"/>
 </g>
 <g transform="translate(0,2424)">
  <path transform="translate(-4) scale(1.8)" d="M18.863,16.496l-7-12C11.685,4.189,11.355,4,11,4s-0.685,0.189-0.863,0.496l-7,12c-0.182,0.311-0.182,0.691-0.004,1.002S3.643,18,4,18h14c0.357,0,0.689-0.191,0.867-0.502S19.044,16.807,18.863,16.496z" fill="#c9c9c9"/>
  <circle transform="translate(-4) scale(1.8)" cx="10.998" cy="14.999" r="1.051"/>
  <polygon transform="translate(-4) scale(1.8)" points="10 8 12 8 11.65 13 10.35 13"/>
 </g>
 <g transform="translate(0,3362)">
  <path d="m11.834 1.3224-1.175-1.1708-4.6584 4.6416-4.6583-4.6416-1.175 1.1708 4.6583 4.6416-4.6583 4.6416 1.175 1.1708 4.6583-4.6416 4.6584 4.6416 1.175-1.1708-4.6584-4.6416 4.6584-4.6416z" fill="#fff"/>
 </g>
 <g transform="translate(0,1056)">
  <rect width="24" height="24" fill="url(#pattern0)"/>
  <defs>
   <pattern id="pattern0" width="1" height="1" patternContentUnits="objectBoundingBox">
    <use transform="scale(.00059952)" xlink:href="#image0"/>
   </pattern>
   <image id="image0" width="1668" height="1668" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABoQAAAaECAYAAADaIXzeAAAACXBIWXMAABcRAAAXEQHKJvM/AAAgAElEQVR42uzdyY+V553o8ZaQWFhCslSSF0iWkJBZICGV9Egt1tydd2y6r+QN0lVa3fcSuh3HiWMTZ3Di4NjEdoidOBhs4inEhbGNMZjRmLEYi6GgCqooajh1zqk6Y51z2L593vJw053gZqiqM7yfxecfOJt6fr9vPc/7D1EU/QMAAAAAAADty48AAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAAAgCPkRAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAQBACAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAYOZUazc7qrXaw9OqtUcq1dr6v9JV1w0AALSXUnnqZKFYOh3LTkzuSI1nXvta/9WBxy5f6fvO5b7+aVe+cfU7V/qvfufgoSP/+P62D5d0ffDRtG3bP572wYexHUu2f/TJwg8/ju1c+NGOTx/4+JNPF3xp131mMAAEIQCY1ejzX2LPdOSZqlRTdREAANB+SuWpKF8oRdnJXDqTnTg3NDzSdX1oeHPv5b51p8/2rDl+8vSqP739XnjrnT+Ht97dOu3tunfe+0t458/vh3fr3tvaFd77y7bw569sff+DsLVre/hL3fvbPgxdH3w0bdv2j6d98GFsR9j+0Sfhw49jO8NHOz4NH3/ytV1hx85d4ZNPd9d9tmTnrs+WfLp7z8JPd++NLdj12d755jcABCEAuL3bPssr1drqr8KP6AMAAG2uPFWJ8oVilJ2YTI+lxo8MXr+x+VzPhbVHjnev2vTGW2Hzm3Vb3p72xp/eCW/G3no3bHn7vdDgIBR27vosfLp7T93eabs+2xt2f7Yv7N6zb+lne/cv2rP3wMI9+w4s2Lv/4DzzHgCCEABJjj8PfRV/Nn0VfwzEAADQ5grF0nT8GR0bP3K5r39D98nTa157/Y0Q++OmN8PGTVvCxs1bwutv/Cm0cBAKn+3dH/bsPRD27DsQ9u4/GFu2b//ni/cd+Hzh/oOHFpgJARCEAEhCAOpy8wcAAJIhvv0zns4ODA7d6Dp95tza3Xv2r3z1tU3h93/cFP6wcXN4beOXMSgBQSjs2/952Hfg87D/4KFpBz7/YsnBzw8vPHjosEAEgCAEQEsHoI6vvvsjAAEAQIK+/ZPJTqaHhkd39Vy4uG5r1/YVv/v9xhB75Q8bw6t/eD0IQt8EoXDw88Ph4KEvff7FkSWHvjjywKHDR+8zUwIgCAHQCreA1noCDgAAknULaCyVHrjUe2XDwUOHV738uz+E377yWtjwauyPQRC67SAUDsUOHw1fHDm27PCRY4sOHz1+v1kTAEEIgKaKQPVBsM8wDAAAyTCZK0Qjo2NHzvZcWPfu1q4VL/721fDShlfDyxt+HwShGQlC4XDs6PFw5OjxzrpFR46dEIcAEIQAEIEAAIDZVSiWopGxVM/Zc+fXvf3eX1b85uXfhd+8/EqIY5AgNKtB6EvHToSjx090HjvevejYiZPiEACCEACzp1Ktra7baxgGAIBkKJamolQ6k7lwqXfDRzs+Xfn8b34bXnhxQ1j/UhyDBKEGBKFw7Hh3OHbiZDh+4uSyE92nHjxx8tR88yqAIAQAM3UbaFN9GKwYiAEAIClPwuWj60PDu744cnTNr9e/HGJxDBKEmioIhRPdp8KJk9OWdp883dF96sw8cyyAIAQAd3MbqNswDAAAyVCeqkSp8Uzm/MXeDVveenfFuhdeDM+98FIQhFoiCIXuk6dD96kznSdPnXnw1Omzbg0BCEIA8K23gToq1dr6+jCYMhADAEAy5IulaHh0rOfo8e61zz63Pvzq178J655/MQhCLRmEwsm6U6fPhlNnzi4+febcArMugCAEAJ6FAwCABMvlC9G1weu7t3348cpfrnsh/PK59UEQaqsgFE6fORdOnz23tK7D7AsgCAEgBHUZhgEAIDmyE5PVK31Xt3V98PHKX/zq+TAdgwShdg5C086c7Vl29tx5YQhAEAJACAIAANo9BF24dHnL65v/tOLnz/46PPPs80EQSlQQCmfPnY8tO9dzQRgCEIQAEIIAAIB2MjGZmw5Bf9y0ZcXPfrEu/PyXzwVBKNFBKJzruRDOnb+wrOf8RWEIQBACoM1CUIcQBAAAyftG0NVrg7u3dm1f+ZNnfhV++sy6IAgJQn8VhELP+Yvh/IWLy+qEIQBBCIA2CEHr68NgxUAMAADJUCyVo4HBoaNb39++8ic/fzbEMUgQEoS+JQh95dKSCxcvLTBLAwhCALSYSrW2uj4MpgzEAACQDOWpSjQyOjaw78Dna378s1+Gp3/2bBCEBKE7CELhwsVY76KLly7PN1cDCEIANP+toOWVaq3bQAwAAMmRyU5WT53peWXtT54Ja3/6iyAICUL3EITCxUuXOy/2Xl5oxgYQhABo3ufhNhmGAQAgOfKFYtR/bWD3q6+9vuKpp58JgpAgNENBKFzsvRwu9V5Z1nv5imfkAAQhAJomBlVrj/hOEAAAJEdpqhINj4wN7N1/cM2TT/88xAQhQWgWglDovTxtce/lvnnmbwBBCIDG3graayAGAIDkmMwXop7zl7Y8sfan4Uc//lkQhAShOQhCdX2dl6/0PWAWBxCEAHArCAAAmM1bQeUvbwV99Mmnq5546qdBEBKE5jgIhctXYv1LrvT1zzeXAwhCALgVBAAAzPStoFwhOnf+4pYfPPl0+OFTPwmCkCDUwCAUrvT1d17pv+q2EIAgBIBbQQAAwEzeCvrw452rHv/R00EQEoSaJAiFK/1XQ1//1cX9V6/5thCAIATADN8K2mQgBgCA5MgXitHF3ivbHn/ix2GaICQINV8QCv1Xr3XWLTC7AwhCANx7DFpeHwb7DMQAAJAc4+lsdfeefWu+/8O1QRAShJo8CH3tQTM8gCAEwF2qVGurPREHAABJeiJuKhq4fqPnpQ2/X/HYD58KgpAg1EJBKFy9NrC0br55HkAQAuDOnojrMhADAECynog723Nhy6OPPxm+94OngiAkCLVgEIp1XhsY9IQcgCAEwG3EoIc8EQcAAMmSzk5UDx46/OSj3/9REIQEoRYPQuHawGBsoRkfQBAC4JYxqPawJ+IAACBZbgyPDmz7cMeq//j+E0EQEoTaKAiFgcHriwcGh+aZ9wEEIQD+6/eC1hqGAQAgWd8L6r86cHT9y6+s+PfHngiCkCDUhkGobmhpne8KAQhCAHwVg3wvCAAAEva9oAsXe7et+d4PQxyDBCFBqI2DUKxz8PrQfeZ/AEEIIMnfC+qoVGvdBmIAAEhWDDp89Pi6NY/+IAhCglBCglAYvD4Url+/0WEXACAIASQyBtWHwT4DMQAAJEc6M1HdueuzNd999PEgCAlCCQxC4frQjQfsBAAEIYAkxaDl9WGwYiAGAIAkxaBs9f0PPlq1+j8eD4KQIJTgIBSGhoYX2Q0ACEIAYhAAANB2rg8ND77+xlsr/9+/fz8IQoKQIDQchm6IQgCCEEA7x6Bq7RExCAAAkheDnlv/0or/u+axIAgJQoLQN0Eo3BgeWVo3z74AQBACaCuVam21YRgAAJIag74XBCFBSBD6myAkCgEIQgBiEAAA0NoGh24MPvfC1zFIEBKEBKFbBKHpKDQ8MioKAQhCAGIQAADQejFo3fMvrvi3734dgwQhQUgQ+pYgFIZHRkUhAEEIQAwCAABaLwb96+pHgyAkCAlCtx2EpqPQyOiYKAQgCAGIQQAAQOvEIEFIEBKE7jgIhZHRMVEIQBACEIMAAIDWiUGCkCAkCN1VEJqOQqNjKVEIQBACaG7V2s3lhmEAABCDBCFBSBC66yAURsdSS+0YAAQhgGaPQRUDMQAAJMfQjZGBvxeDBCFBSBC6pyAUW2TXACAIAYhBAABAw6Uz2erWru2r/l4MEoQEIUHonoNQGEuJQgCCEEBzxaCO+jDYZyAGAAAxSBAShAShGQ1CsYV2DwCCEIAYBAAAzLlcoRjtP3DoyW+LQYKQICQIzVgQqhvvsIMAEIQAGqpSrXUZiAEAIFkx6NDhY+v+pxgkCAlCgtCMBqGQGh+/zx4CQBACaFQM2mQgBgCA5CiVp6KLly7vuZ0YJAgJQoLQjAehztR4er59BIAgBDDXMWi1gRgAAJKl/9rgkduNQYKQICQIzXgQqksvHU+n59lLAAhCAHP13aDl9WGwYiAGAIDkGLoxMrDu+RdXCEKCkCDU0CAUxtPpxXYTAIIQwFzEoI76MJgyEAMAQHKkM9nq1q7tq+4kBglCgpAgNGtBqC6z0I4CQBACmO2n4roNxAAAkBy5QjHaf+DQk3cagwQhQUgQmtUgFNKZzP32FACCEMBsxaD1BmIAAEiOUnkq6rlwadvdxCBBSBAShGY9CHWmM9n59hWAIORHAJjhp+JqDxuIAQAgWQaHbgzebQwShAQhQWjWg1BddqmdBSAI+REAZvq7QRUDMQAAJOu7QRs3b1kpCAlCglBTB6HYg3YXgCAEgO8GAQAAc/rdIEFIEBKE5jwIhUw263tCgCAEgO8GAQAAd+ZevhskCAlCglBDglBnJjsxzx4DEIQAuNun4pYbhgEAIFmGbowMrHv+xRWCkCAkCLVUEKqbWGyXAQhCANztd4P6DMQAAJAck7l8tLVr+6qZiEGCkCAkCM15EArZ7MQDdhqAIATAnT4Vt8lADAAAyVEqT0WnzvRsmakYJAgJQoJQQ4JQZ3Zicr69BiAIAXCbt4NqDxuIAQAgeU/FzWQMEoQEIUGoIUEoZCcml9htAIIQALelPgymDMQAAOCpOEFIEBKEWjIIhYmJSU/HAYIQAP/jU3HrDcQAAOCpOEFIEBKEWjoIdU5M5jwdBwhCANzqqbibyw3EAACQLCOjqcxsxCBBSBAShBoahMLEZG6xXQcgCAFwq9tB3QZiAABIjlyhGO3YuWuNICQICUJtGYTC5GTufvsOQBAC4L/HoNUGYgAASJbeK/27ZysGCUKCkCDUFEFoWd08ew9AEALg66fiOurDYMVADAAAyZHOZKvrnn9xhSAkCAlCbR2EYgvtPgBBCICvbwdtMhADAEBylMpT0YmTpzfMZgwShAQhQahpglCYzOXm238AghCA20EPGYgBACBZRkZTmdmOQYKQICQINVUQWmwHAghCAG4HdRuIAQAgOYqlcrRj5641gpAgJAglKgiFXC6/wB4EEIQAEns7qPawgRgAAJJlcOhGz1zEIEFIEBKEmi4ILbULAQQhgISqD4N9BmIAAEiOyVw+2tq1fZUgJAgJQokMQiGXz3fYhwCCEEDynopbbSAGAIBk6b3Sv3uuYpAgJAgJQk0ZhJbZiQCCEEDybgelDMQAAJCs20EbN29ZKQgJQoJQooNQyOcLbgkBghCA20EAAIDbQYKQICQItXkQ6swXCvPsRwBBCMDtIAAAwO0gQUgQEoTaNwiFfKGw0H4EEIQA3A4CAADcDhKEBCFBqL2DUGehUHRLCBCEANwOAgAA3A4ShAQhQaiNg1AoFIoP2JMAghCA20EAAIDbQYKQICQItXcQWmZXAghCAG4HAQAAbgcJQoKQINTeQSgUisUO+xJAEAJoM9Vq7REDMQAAJEtf/7VdjYpBgpAgJAi1RBBySwgQhADa8Lm4bgMxAAAkR7FUjnbs3LVGEBKEBCFB6FuCUOx+exNAEAJol9tBtZvLDcQAAJAsg0M3ehoZgwQhQUgQapkgtMTuBBCEANrndlCXgRgAAJKjVJ6KDh0+tk4QEoQEIUHoNoJQKBZL8+1PAEEIoPVvB3UYiAEAIFlS4+l0o2OQICQICUItFYQW2aEAghBA698OWm8gBgCAZDl1pmeLICQICUKC0B0Eoc66efYogCAE0MLqw2DKQAwAAMkxmctHGzdvWSkICUKCkCB0B0Eo1mGPAghCAK36XFy19oiBGAAAkuXa4NCRZohBgpAgJAi1XBBaapcCCEIArftcXJeBGAAAkqNUnor27D2wVhAShAQhQeguglAolkr32acAghBAq90Oqt3sMBADAECypMbT6WaJQYKQICQItWQQWmSnAghCAK13O2itgRgAAJKl58KlbYKQICQICUL3EIQ67VQAQQigxdSHwT4DMQAAJEexVI62dm1fJQgJQoKQIHQPQSiUSuX77VUAQQigdZ6Le8hADAAAyTJ0Y2SgmWKQICQICUItG4QW260AghCA5+IAAIAmdeLk6Q2CkCAkCAlCMxCEQqlcnme/AghCAK3xXFzKQAwAAMmRKxSjjZu3rBSEBCFBSBCaoSDUYb8CCEIAnosDAAA8FycICUKCUHsHIc/GAYIQgOfiAAAAz8UJQoKQINTmQSiUy1OejQMEIYAmfy6uz0AMAACeixOEBCFBSBC6xyDk2ThAEALwXBwAANAsUuPpdDPGIEFIEBKEWj4ILbJrAQQhgOZ9Lm61gRgAAJKl58KlbYKQICQICUKzEIQ67VoAQQigeYPQXgMxAAAkR6k8Fe3YuWuNICQICUKC0CwEoVCemlpg3wIIQgDN+f0gQzEAACRIOpOtNmsMEoQEIUGoLYLQQvsWQBACaLrvB9UeNhADAECyXBscOiIICUKCkCA0i0FoqZ0LIAgBNN9zcZsMxAAAkCwnTp7eIAgJQoKQIDSLQSg2z94FEIQAmuu5uD4DMQAAJEeuUIw2bt6yUhAShAQhQWiWg9D99i6AIATQNM/F3ewwEAMAQLKkxtPpZo5BgpAgJAi1TRB60O4FEIQAmiUIVWuPGIgBACBZ+vqv7RKEBCFBSBCagyDkO0KAIATQRN8PWm8gBgAA3w8ShAQhQUgQmoUgFKZ8RwgQhACaJgh1G4gBACA5iqVytLVr+ypBSBAShAShOQpCviMECEIAzcBADAAAyZLOZKvNHoMEIUFIEGqrILTQ/gUQhAAa/f2g2s3lBmIAAEiWoRsj5wQhQUgQEoTmMAgtsYMBBCGAxj8Xt9ZADAAAyXL+Yu9mQUgQEoQEoTkMQp12MIAgBND4INRlIAYAgGTZs/fAWkFIEBKEBKE5DEJ1lfn2MIAgBNDYINRtIAYAgOTIFYrRxs1bVgpCgpAgJAjNcRC63x4GEIQAGshADAAAyZLOZKutEIMEIUFIEGq7ILTQHgYQhAAapFq7udxADAAAyTI8MnZOEBKEBCFBqAFBaIldDCAIATQqCFVrjxiIAQAgWS719nUJQoKQICQINSAILbOLAQQhgMZ9P2i9gRgAAJLlxMnTGwQhQUgQEoQaEISCXQwgCAE0LgjtNRADAECy7Ni5a40gJAgJQoJQI4LQVKWywD4GEIQAGhOEug3EAACQHJO5fLTu+RdXCEKCkCAkCDUoCN1vHwMIQgANYCAGAIBkyU5MRq0SgwQhQUgQassgtNA+BhCEAOZYtXazw0AMAADJMjwydk4QEoQEIUGogUFokZ0MIAgBzHkQqj1sIAYAgGQZujEiCAlCgpAg1MggtMROBhCEAOY6CFVrjxiIAQAgWc5f7N0sCAlCgpAg1MAgtMxOBhCEAOZYpVpbbyAGAABBSBAShAQhQWgOg1CwkwEEIQBBCAAAmGV79h5YKwgJQoKQINTIIFSpVOfZywCCEMDcBqFuAzEAACTLjp271ghCgpAgJAg1OAgtsJcBBCEAQQgAAJglxVI52tq1fZUgJAgJQoKQIAQgCAEJUh8I+wzFAACQHJO5fNRKMUgQEoQEobYNQh32MoAgBDC3QchQDAAAgpAgJAgJQoLQXAehhfYygCAEIAgBAACzJJ3JVgUhQUgQEoQEIQBBCBCEAACANjY8MnZOEBKEBCFBqAmC0IP2MoAgBDBHqrWbDxmIAQBAEBKEBCFBSBBqQBBaYjcDCEIAcxaEag8biAEAQBAShAQhQUgQEoQAQciPAAhCAACAICQICUKCkCAkCAGCEIAgBAAAtIpLvX1dgpAgJAgJQoIQgCAECEIAAEAbO3+xd7MgJAgJQoKQIAQgCAGCEAAAIAgJQoKQICQICUKAIAQgCAEAAIKQICQICUKC0D0FoU67GUAQAhCEAAAAQUgQEoQEofYOQsFuBhCEAAQhAABAEBKEBCFBSBACEIQABKHWVZ6qRIViKcpO5AEAEiNfKEWl8pTzYBOoVGvrzUMAAIIQIAgxS3L5YpQaz0bDI+MAAIk1lspOn4ucDwUhAABBCEAQaivFUnl68WEBBADw/42OZaZvTTsvCkIAAIIQgCDUFreCLHwAAG7NbSFBCABAEAIQhMQgAIAEiL8x5PwoCAEACEIAglDLiZ8/sdwBALh9+YLn4wQhAABBCEAQaiHlqcr0m/gWOwAAt29kND19jnKeFIQAAAQhAEGoJcRPnljqAADcuXRm0nlSEAIAEIQABKHWEP93q4UOAIBbQoIQAIAgBCAItan47XvLHACAu5fLF50rBSEAAEEIQBDyXBwAgGfjEIQAAAQhAEGogVLjWYscAIB7EJ+nnCsFIQAAQQhAEBKEAADa2OhYxrlSEAIAEIQABCFBCACg3TlXCkIAAIIQgCAkCAEAeDIOQQgAQBACEIQaJ/4IskUOAIAgJAgBAAhCAIJQG8vlixY5AAD3IDuRd64UhAAABCEAQai5lcpTFjkAAPegWCo7VwpCAACCEIAg1PzG0xOWOQAAnosThAAABCEAQaidFYolCx0AgLsQn6OcJwUhAABBCEAQahmZbM5SBwDgDsS3rJ0jBSEAAEEIQBBqOWOprOUOAMBtiM9N5amKM6QgBAAgCAEIQq0nXmqIQgAAYpAgBAAgCAEIQgmIQunMpGUPAMAtnokTgwQhAABBCEAQahvxB5JT424LAQDERscyUb5Qck4UhAAABCEAQag9FUvlKJPNTcehkdG0hRAAkBjx+Sc+B8X/KONcKAgBAAhCAIIQAAAgCAEACEIAghAAACAIAQAIQgCCEAAAIAgBAAhCAIIQAAAIQgAACEKAIAQAAAhCAACCEIAgBAAACEIAAIIQgCAEAAAIQgAAghCAIAQAAAhCAACCEIAgBAAACEIAAIIQgCAEAAAIQgAAghCAIAQAAIKQIAQAIAgBghAAACAIAQAIQgCCEAAAIAgBAAhCAIIQAAAgCAEACEIAghAAACAIAQAIQgCCEAAAIAgBAAhCAIIQAAAgCAEACEIAghAAACAIAQAIQoAgZCgGAABBCABAEAIQhAAAAEEIAEAQAhCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAAEEIAEAQAhCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAQBACAEAQAgQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIUAQEoQAAEAQAgAQhPwIgCAEAAAIQgAAghCAIAQAAAhCAACCEIAgBAAACEIAAIIQgCAEAAAIQgAAghCAIAQAAAhCAACCEIAgBAAACEIAAIIQgCAEAACCkHkIAEAQAgQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQAQYi5U56qRIViKZrMFaLsRB4AaAPx3/b4b7yzDoIQAIAgBCAIJVy+UIrG0xPR8Mg4ANCm4r/1uXzR2QdBCABAEAIQhJKmWCpHqfGsJRkAJMhYKjt9BnAWQhACABCEAAShBIj/Q3hkNG0xBgAJ5bYQghAAgCAEIAglIAZZhAEAohCCEACAIAQgCLXxM3EWYADA1wrFks6ZO3MAACAASURBVDMSghAAgCAEIAi1k/JUJRody1h+AQDfiM8G8RnBWQlBCABAEAIQhNpEdiJv8QUA/I34jOCshCAEACAIAQhCbcLtIADg7xkZTTsrIQgBAAhCAIJQO4i/D2DhBQDcSr7gW0IIQgAAghCAIOS5OACgrWWyOWcmBCEAAEEIQBBqdanxrGUXAHBL8VnBmQlBCABAEAIQhAQhAEAQAkEIAEAQAhCEBCEAQBACQQgAQBACEIQEIQBAEAJBCABAEAIQhGZHOjNp2QUA3NJ4esKZCUEIAEAQAhCEWl0uX7TsAgBuaTJXcGZCEAIAEIQABKFWVypPWXYBALcUnxWcmRCEAAAEIQBBqA3ET8FYeAEAvh+EIAQAIAgBCEJtrFAsWXoBAH8jPiM4KyEIAQAIQgCCUBvJZHMWXwDAN+IbxM5ICEIAAIIQgCDUZspTlWgslbUAAwCmzwTx2cAZCUEIAEAQAhCERCEAQAwCQQgAQBACEIRaNQrFT8RYiAFAMp+JE4MQhAAABCEAQShB8oVSNDqWsRwDgASI/+bHf/udgRCEAAAEIQBBKKEKxVKUyeai1Lin5ACgncR/2+O/8fHfemceBCEAAEEIQBACAAAEIQAAQQhAEAIAAAQhAABBCEAQAgAABCEAAEEIQBACAAAEIQAAQQhAEAIAAEEIAABBCBCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAAEEIAEAQAhCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAAEEIAEAQAhCEAABAEBKEAAAEIUAQAgAABCEAAEEIQBACAAAEIQAAQQhAEAIAAAQhAABBCEAQAgAABCEAAEEIQBACAAAEIQAAQQhAEAIAAAQhAABBCEAQAgAABCEAAEEIEIQAAABBCABAEAIQhAAAAEEIAEAQAhCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAAEEIAEAQAhCEAAAAQQgAQBACEIQAAABBCABAEAIQhAAAQBACAEAQAgQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIUAQMhADAIAgBAAgCPkRAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAEITMRAIAgBAhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCzaZQLEW5fDHKTuQBANreZK4wff4pT1WcBQUhAABBCEAQav8INJ6eiIZHxgEAEis+D8X/GON8KAgBAAhCAIJQWymVp6LUeNYCCADgr4ylslGxVHZeFIQAAAQhAEGo9cX//Toymrb0AQC4BbeFBCEAAEEIQBBq+RhkyQMAIAoJQgAAghCAINSm4udPLHcAAG5fvlByjhSEAAAEIQBBqLWMjmUsdgAA7kD8zG55quIsKQgBAAhCAIJQa8hO5C11AADuQnyOcp4UhAAABCEAQcjtIAAAt4QQhAAABCEAQaixCsWSZQ4AwD3I5YvOlYIQAIAgBCAIeS4OAKCdpTOTzpWCEACAIAQgCDW31HjWIgcA4B7E5ynnSkEIAEAQAhCEBCEAgDY2lhKEBCEAAEEIQBAShAAA2p5zpSAEACAIAQhCghAAgCfjEIQAAAQhAEGoceKPIFvkAAAIQoIQAIAgBCAItbHJXMEiBwDgHmQn8s6VghAAgCAEIAg1t1J5yiIHAOAeFEtl50pBCABAEAIQhHxHCACgXY2OZZwnBSEAAEEIQBBqDYViyUIHAOAu5Asl50lBCABAEAIQhFpHJpuz1AEAuAPxLWvnSEEIAEAQAhCEWkp5qhKNpTwdBwBwu0/Fxecn50hBCABAEAIQhEQhAIA2NDKajoqlsvOjIAQAIAgBCEKtHYXG0xOWPQAAt3gmzs0gQQgAQBACEITaRvyB5PgpFIsfAIAvn4jL5YvOiYIQAIAgBCAItW8YSmcmPSUHACROfP6Jz0Hxeci5UBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAAAQhAAAEIQAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAAAQhQQgAQBACBCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhAAEIQAAQBACABCEAAQhAABAEAIAEIQABCEAAEAQAgAQhABByFAMAACCEACAIAQgCAEAAIIQAIAgBCAIAQAAghAAgCAEIAgBAACCEACAIAQgCAEAAIIQAIAgBCAIAQAAghAAgCAEIAgBAACCEACAIAQgCAEAgCAEAIAgBAhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCAACAIAQAIAgBghAAACAIAQAIQgCCEAAAIAgBAAhCAIIQAAAgCAEACEIAghAAACAIAQAIQgCCEAAAIAgBAAhCAIIQAAAgCAEACEIAghAAACAIAQAIQoAgJAgBAIAgBAAgCPkRAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAQhAAABCEAQQgAABCEAAAEIQBBCAAAEIQAAAQhAEEIAAAEIfMQAIAgBAhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCAACAIAQAIAgBCEIAAIAgBAAgCAEIQgAAgCAEACAIAQhCAACAIAQAIAgBghBzq1AsRflCKcpO5AEAZtRkrjB91iiVp5y7EIQAAAQhAEGoEREonZmMRkbT0fDIOADArBsdy0xHovJUxXkMQQgAQBACBCFmU/zfuanxrKUUANAw8T+kxGHI2QxBCABAEAIEIWZB/CycG0EAQLOI/0nFbSEEIQAAQQgQhJhBuXzR4gkAaDpjKVFIEBKEAAAEIUAQYkYUS2U3gwCApr4p5MwmCAEAIAgBghD3KP7PW8smAKCZTeYKzm2CEAAAghAgCOGpOACgncW3mT0dJwgBACAIAYIQd2l0LGPJBAC4JYQgBAAgCAEIQu387SDLJQCgVcTP3DrDCUIAAAhCgCDEHcpO5C2XAICW4tk4QQgAAEEIEIS4Q+PpCYslAKClFIol5zhBCABAEPIjAIIQdyI1nrVYAgAEIQQhmso//7bWF/unb1S/9PJ/V+n7P69Vt//LxuqbX/vum9WnH3u7+r9jP3in+r/8ngAIQvCf7N1LjN3XfdhxwGCBLNlstFXbRVc1tAwqW6bcNrbRJBVsN5JjB2VbRXVrO2Xc1k89aFmp7ViyJNrmvDj0NG1dt2lQARbfgaAuGiCwFyxatFoUMTVz3+87I5uMsrid/yWHHIkzw5m5/8f5n/9n8VkIFkB55p7De3/fe84fBCEEIQBAEEIQIkAf/P23JlPPbUwefof1d/r6eAejO54dTY5NDSd//1ujwT98cfzGJ06Nf/I7i+srj2/6/B9uPPbp5Y2P+pkDIAgBCEKCEACAIIQgRARB6J0GN33tjr/3+8PrH//O6I1PfW/02uML45Xf+3fjx77wH9ff6/cBgCAEIAhFodnqGiwBAIIQghCVD0J39G/7wMlEb/KxFwZvfPK7w9eeWBy9eGJl/JjfEQCCEIAgVDrd3sBgCQAoFe/hBCEEobyD0N26k498o9//rVOD155YGL74xOLItXMACEIAglDYRuN1gyUAoDQazY73cIIQglAQQei2ZxKdqY8+33vjn5werPzOwuiJzf/+o36XAAhCAIKQ5wgBABxCf+C6OEEIQSjcIHRHe/KBp9uTX/tmb/WTp/r/9fH5oUAEgCAEIAgVL7mH34AJAAhdrd723k0QQhAqVRB66B1ak0f+oPt/Hp/rv3jiB4O/4/cMgCAEIAgVIrl+xaAJAAhZ8iUW79sEIQShMgeh7T78XHvw6Iu9K/98qf8Zv3MABCEAQSg34/WN6bduDZsAgBB1ewPv2QQhn4kEoaiC0ENPJZo3bf7zx57v/tkT872n/80fDu7zGgBAEAIEIUFIFAIAKqfZ6nqvJggJQoJQ3EHotsbk/Zs+/nz7JzfjUF8cAkAQAgQhsotC9YYoBAAUb3WtOen1h96jIQgJQrtHoUiD0NSTifrko9/u/Nk//n7vy5s/j6NeGwAIQoAgROqS4ctarWUYBQAUdipoNF73vgxBSBCqfBDa8sFnGtcf/U77tU9+d3DcawQAQQgQhEhdfzCaDmTEIQAga8kp5XanLwQhCCEI7RCE7qhNPvT1xuCTL3fO/Pb3hn/T6wVAEAIQhAAAAEEIQSjCIDT11Zs+9u3mTz55qv+vvW4ABCEAQQgAABCEEIQiDULv/+ra1K8+W5+eGvrUd50aAhCEAAQhAABAEEIQijII3bb5v/3mC83XPvHy4Ne8lgAEIQBBCAAAEIQQhCIMQu/b8pW1yW98o/7Gb73cc50cgCAEIAgBAACCEIJQrEHofV9ZnfrVr9UG//T77ac3f6ZHvb4ABCEAQQgAABCEEIQiDEJbHn66dv3R73TmT5zt3Od1BiAIAQhCAABAMMaCkCAkCKUWhG56c/LwU6vXP/VSY0UYAhCEAAQhAAAgiBg0XheEBCFBKO0gtOVOGGoLQwCCEIAgBAAAFBeDBCFBaO8gtC4IzRCE3vflxLXbYcgzhgAEIQBBCAAAKCQG3QxCbwlCgpAglGEQ2nLsqdXrv/lCe14YAhCEAAQhAAAg1xg0Xt8QhAQhQSinIPTgLX/3mTcHv/1y68teiwCCEIAgBAAA5BKDBCFBSBDaJQg9mV0QevBLP5v68LNrq0/MNR/zmgQQhAAEIQAAINMYJAgJQoJQcUFoy0eea17d/H3c77UJIAgBCEIAAEAmMUgQEoQEoeKDUPLn3PqdvOT5QgCCEIAgBAAApB6DBCFBSBAKKgglRpuOe50CCEIAghAAAJBaDBKEBCFBKLggtOX1TQ94vQIIQgCCEAAAMHMMEoQEIUEo2CC05aRr5AAEIQBBCAAAmCkGCUKCkCAUfBBKXNt0zGsXQBACEIQAAIBDxSBBSBAShEoRhLasOC0EIAgBCEIAACAGHTgGCUKCkCBUqiCUGG16xOsYQBACEIQAAEAM2ncMEoQEIUGodEFoyytOCwEIQgCCEAAAiEGCEIJQ3EFo67SQZwsBCEIAghAAAIhBghB3+9A337q+FYQ+KAiVOQhteclpIQBBCEAQAgAAMUgQ4h0ePfXzNwShqIJQ4uqmB7y+AQQhAEEIAADEIEEIQSjeILTlhNc4gCAEIAgBAIAYJAghCN0OQo0Yg1DiFVfIAQhCAIIQAACIQYKQICQIxR2EEtdcIQcgCAEIQgAAIAYJQoKQIBR3EHKFHIAgBCAIAQCAGCQICUKCUEWCUGLFFXIAghCAIAQAABWOQYl1QUgQOmwQ+rogVJIglLjqCjkAQQhAEAIAgIrGIEFIEBKEKhOEEqNNj1gDAIIQgCAEAAAVi0GCkCAkCFUqCHmuEIAgBCAIAQBAFWPQNAhtCEKCkCBUsSDkuUIAghAgCAlCAABQpRgkCAlC5QhC3fCC0FdLH4S2niskCgEIQoAgBAAAxB6DBCFBSBCqdBBKXNv0gHUBIAgBghAAABBxDBKEBCFBqPJBKDHadMzaABCEAEEIAACINAYJQoKQICQIbXPc+gAQhABBCAAAiDAGCUKCkCAkCIlCAIIQIAgBAACRxyBBSBAShAShHaxYJwCCECAIAQAAEcUgQUgQEoQEIVEIQBACBCEAACDyGCQICUKCkCAkCgEIQoAgBAAARB6DBCFBSBAShO7h6qaj1g0gCAEIQgAAQIljkCAkCAlCgpAoBCAIAYIQAAAQeQwShAQhQaj4IJT8u4EHIVEIEIQABCEAAKDMMUgQEoTKGYQ6UQWhB7/052UIQqIQIAgBCEIAAEBZY5AgJAgJQoKQKAQgCAGCEAAAEHkMEoQEIUFIEBKFAAQhQBACAAAij0GCkCAkCAlCohCAIAQIQgAAQOQxSBAShAQhQUgUAhCEAEEIAACIPAYJQoKQICQIzWjFmgIEIQBBCAAAxKDAY5AgJAgJQiEEoZ+VOQiJQoAgBCAIAQCAGCQIUekg9Gx4QeghQUgUAhCEAAQhAACoWgwShAQhQUgQStEJ6wsQhAAEIQAAEIMEIQQhQSjuIJQ4bo0BghCAIAQAAGKQIIQgJAjFHYQSj1hngCAEIAixi+FoPBkMR5NubzBpd/oAAKnpD0bT9xm3Bv+IQYIQMwahsSAkCN3LaNMD1hogCAEIQtySDGaare5kda05eXO1AQCQuVq9Pf0CijgkBglCgpAgJAjlEIWOWm+AIAQgCFXaaLw+aTQ7hlIAQGGSL6QkYch7MzFIEBKEBCFBKENXRSFAEAIQhCp9KsiJIAAgFMmXVJwWqnYMEoQEIUFIEMrYijUHCEIAglDlJPf3GzwBACFeIycKVTcGCUKCkCAkCOXgpHUHCEIAglBlDEdjJ4MAgKBPCnnPVs0YJAgJQoKQIJST49YeIAgBCEKVkHzz1rAJAAiZZwpVMwYJQoKQICQI5WS06QHrDxCEAAShqPX6Q0MmACB4yWlmV8dVLwYJQoKQICQI5ejapqPWICAIAQhC0VqrtQyZAACnhMQgQQhBSBCqehBKvGINAoIQgCAU7bODDJcAgLJIrrn1Hq5aMUgQEoQEIUGoACetQ0AQAhCEotPu9A2XAIBScW1ctWKQIFRNn17+xUpaQehhQUgQOpxj1iIgCAEIQlFpNDsGSwBAqQyGIzGoQjFIEBKEBCFBqCAjzxMCBCEAQSgq9UbbYAkAEITEIEEIQUgQEoTu9rr1CAhCAIKQIAQAIAiJQYIQglDgQWhNEPI8IUAQAhCEEIQAAEFIDBKEEIQEIUHI84QAQQhAEKqEZqtrsAQACEJikCCEICQICUK7u+Z5QoAgBCAIlV63NzBYAgBKRQwShBCEBCFBqACvWJuAIAQgCJXaaLxusAQAlEaj2RGDBCEEodyC0M0oFFoQqgtCxXnE+gQEIQBByHOEAABy0OsPxSBBCEFIEBKEijJydRwgCAEIQqWW3MNvwAQAhG6t1hKDBCEEIUFIECra69YoIAgBCEKllly/YtAEAIQs+RKLGCQIIQgJQoJQAE5Yp4AgBCAIlXf4sPlBu1Z3dRwAEKZ2py8GCUI+EwlCgpAgFNLVcfdbq4AgBCAIldZwNJ5exWLoBACEpNnqikGCkCAkCAlCgpCr4wAEIUAQIu2TQvWGk0IAQBi6vYEYhCAkCAlCglCoHrFeAUEIQBAqvV5/OFldaxpEAQCFSL6gkpxeFoMQhASh0gahZwShilwdd9SaBQQhAEEomjDUaHZcJQcAZC55nmGr3atECBKDBCEEIUEoGivWLCAIAQhCAAAgBglCCEKCUPyOWbeAIAQgCAEAgBgkCCEICUJxu2bdAoIQgCAEAABikCCEIJRhEKoJQmE4ae0CghCAIAQAAGKQIIQgJAjFbbTpfusXEIQABCEAAMQgMUgQQhAqbxBKfheiz72sWL+AIAQgCAEAIAaJQYIQglBpg1DycxN89uWYNQwIQgCCEAAAYhCCEIKQIBS3q9YwIAgBCEIAAIhBCEIIQoJQ/I5bx4AgBCAIAQAgBiEIIQgJQnG7tumotQwIQgCCEAAAYhCCEJULQu3wgtBXBKEMnbSWAUEIQBACAEAMQhBCEBKE4jZySggQhAAEIQAAxCAEIQQhQSh+L1nPgCAEIAgBACAGIQghCAlC8bvfmgYEIQBBCAAAMQhBCEEo1SD0fkEoNCvWNCAIAQhCAACIQQhCCEKCkFNCAIIQgCAEAIAYhCAkCAlCgpBTQgCCECAIAQCAGCQIIQgJQoKQU0KAIAQgCAEAgBgkCCEI7TcIDQQhQcgpIUAQAhCEAAAQg8QgQQhBSBDCKSFAEAIQhAAAEIMQhBCEBCGcEgIEIQBBCAAAMQhBiDyD0Ci8IPR0eEHofYKQU0KAIAQgCAEAIAaJQYIQgpAgxMxessYBQQhAEAIAQAxCEEIQEoTiNtp01DoHBCEAQQgAADEIQUgQEoQEobidtM4BQQhAEAIAQAxCEBKEBCFBKG7XrHNAEAIQhAAAEIMQhAQhQUgQit9xax0QhAAEIQAAxCAEoUr7/H+4/hlBSBCK3FVrHRCEAAQhAADEIAShSvvCD68/Fk4Q6gtCglBWjlnvgCAEIAgBACAGIQgJQoKQIBS3FesdEIQABCEAAMQgBCFBSBAShOJ31JoHBCEAQQgAADEIQUgQEoQEobidsOYBQQhAEAIAQAxCEBKEMglCQ0FIEArFNWseEIQABCEAAMQgBCFBSBAShOJ3zLoHBCEAQQgAADGo0kaCkCAkCAlC8Vux7gFBCEAQAgBADKp0DBKEBKEyB6EPBBmEVgWhMB219gFBCEAQAgBADKpsDBKEBCFBSBCqiOPWPiAIAQhCAACIQZWNQaOxICQICUKCUCVctfYBQQhAEAIAQAyqbAwShAQhQUgQqpD7rX9AEAIQhAAAEIMqGYMEoYoHoVtRSBAShCriJesfEIQABCEAAMSgSsYgQUgQEoQEoQq5Zv0DghCAIAQAgBhUyRgkCAlCgpAgVDEP2AMAQQhAEAIAQAyqXAwShAShygahpwQh18YBCEKAIGTQAQCAGFSRGHQzCG0IQoKQICQIuTYOQBACBCEAABCDYo1Bo/G6ICQICUKCkGvjAAQhQBACAAAxKOYYJAgJQoKQIOTaOABBCBCEAABADIo8BglCgpAglHUQelMQcm0cIAgBCEIAAIhBFBuDBCFBSBAShFwbByAIAYIQAABikBgUeQwShAQhQSiMIJT8fxFpcnXCXgAIQoAgZPgBACAGiUGViUGCkCAkCAlCFXXVXgAIQoAgZAACACAGiUGViUGCkCAUfBA6KQiRmaP2A0AQAgQhAADEIDGoEjFIEBKEBCFBqMKO2w8AQQgQhAAAEIMEl0rEIEFIEBKEBKEKW7EfAIIQIAgBACAGUYkYlBgLQoKQICQIVdPIfgAIQoAgBACAGEQlYpAgJAgJQoJQxT1gTwAEIUAQAgBADCL6GCQICUKCkCBUcSfsCYAgBAhC5Cr5ID4YjgAActNPDIozGI5FngBi0DQIrQtCgpAgJAhV1iv2BEAQAgQhcolAzVZ3slZrTd5cbQAAVM7qWnP6figJRKJPMTFIEBKE4g5CLUGIe7InAIIQIAiR3dUsmx/kk8GHIRAAwB31RnsyHDk1lHcMEoQEIUFIEOKtY/YFQBACBCFSlww5km/CGvoAAOx8YqjXHwpBOcYgQUgQEoQEId46aV8ABCFAEEIMAgAoQLc3EINyikGCkCAkCAlCeI4QIAgBghBiEABAYQbDsRiUQwwShAShPYPQc4KQIFQJI/sCIAgBghCpqdXbBjsAAAewVmttxQoxKMMYJAgJQoKQIMTUA/YGQBACBCFmltyDb6gDAHBw7U5PDMo4BglCgpAgJAgxddzeAAhCgCDEzJJvtxroAAAcXHLlrhiUbQwShAQhQUgQYmrF3gAIQoAgxMzPDjLMAQA4vOS0tRiUXQwShAQhQUgQYuqqvQEQhABBiJm0O32DHACAGbTaPTEowxgkCAlCgpAgxE32BkAQAgQhZtJodgxyAABmUG+0xaAMY5AgJAgJQoIQtx2zPwCCECAIcWjJAMMgBwDg8Gr1lhgkCCEIpRSEmoIQezlhfwAEIUAQQhACACiQGCQIka4n/8v19wpCghB3WbE/AIIQIAghCAEAuDIuyhgkCFWXICQIcZer9gZAEAIEIQ6t2eoa5AAACELBxiBBSBAShAQh7rA3AIIQIAhxaN3ewCAHAGAG7U5PDBKEEIQEIfLygP0BEIQAQYhDST5gG+QAABzeYDgWgwQhBCFBiLw8Yn8ABCFAEMJzhAAAcrZWa4lBghCCkCBEnk7aHwBBCBCEOLTBcGSgAwBwCMn1u2KQIEQVg1BPEKIor9gfAEEIEISYSaPZMdQBADiA5JS1GCQIIQgJQuTsdfsDIAgBghAzSYYCyZUnhjsAAPe2utacDEdjMUgQQhAShMid/QEQhABBiJklQ41kuGHIAwCwdwwaDMUgQQhBSBCiMEftEYAgBAhCpHJSqFZvG/YAAOygVm+JQYIQgpAgRNGO2SMAQQgQhEhN8oBkp4UAAO6cCmp3ep4ZJAghCAlChOC4PQIQhABBiNRPC/X6w0mj2RGHAIBKSt4HJV+UuRUlxCBBCEFIECIEJ+0RgCAECEJkbjAcAQAV108M4lbm+BNbDBKEBCFBSBDiLiv2CEAQAgQhAACyPUE8PUW83QZikCCEICQIka/X7RGAIAQIQgAAiEFEFYMEIUFIEBKEuMs1ewQgCAGCEAAAYhBRxSBBSBAShAQh7maPAAQhQBACAEAMEoOiikGCkCB0dxDaEIQEIUHIHgEIQoAgBACAGCQGxRSDBCFBSBAShNjRMfsE4IcACEIAAIhBYlA0MUgQEoQEIUEIQQgQhABBCAAAMYjIY5AgJAgJQoIQO3rEPgH4IQCCEAAAYpAYFE0MEoQEIUEojCD00OafK8IE5aR9AvBDAAQhAADEIDEomhgkCAlCglAYQSj5c0QYQQgQhAAEIQAAMQgxSBBCEBKEEIQAQQhAEAIAEIMQgwQhBKFSBKEdopAgFJzX7ROAHwIgCAEAIAaJQdHEIEFIEBKEiTegLwAAIABJREFUBCEEIUAQAgQhAADEIDEo8hgkCAlCgpAghCAECEKAIAQAgBgkBkUegwQhQUgQEoQQhABBCBCEAAAQg8SgyGOQICQI3TsIrQtCglAVjewTgB8CIAgBACAGiUGCEIKQICQIRc4+AfghAIIQAABikBgkCCEICUKCkCAECEIAghAAgBgkBolBghCCUOmD0JOCkCAECEIAghAAAGKQGCQIIQgJQoKQIAQIQgCCEACAGIQYJAghCAlCgpAgBAhCAIIQAIAYhBgkCCEICUKCkCAECEIAghAAgBiEGCQIIQgJQghCgCAEIAgBAIhBiEGCEIKQIIQgBAhCAIIQAIAYJAaJQYIQgpAghCAECEIAghAAgBgkBglCCEKCkCCEIAQIQoAgBAAgBolBYpAghCAkCAlCghAgCAEIQgAAYhBikCCEICQICUKCECAIAQhCAABiEGKQIIQgJAgJQiVw1F4BghCAIAQAIAYhBglClNqvP//WYCsIfVAQEoTYyTF7BQhCAIIQAIAYhBgkCFFqj576+RuCkCCEIAQIQoAgBAAgBolBYpAghCAkCAlCghAgCAEIQgAAYhBikCCEIFT2INQQhBCEAEEIEIQAAMQgwUUMEoQQhAQhQUgQAgQhAEEIAEAMQgwShBCEBCFBSBACBCEAQQgAQAxCDBKEEIQEIUFIEAIEIQBBCABADEIMEoQoZxD6uiAkCAlCgCAEIAgBAIhBiEGCEIKQICQICUKAIAQgCAEAiEGIQYIQgpAgJAgJQoAgBCAIAQCIQWKQGCQIIQiFF4S+KggJQoAgBCAIAQCIQYhBghCCUIpBqCsIIQgBghCAIAQAIAaJQQhCCEKCEIIQIAgBCEIAgBgkBolBCEIIQoIQghAgCAEIQgCAGIQYJAghCAlCghCCECAIAYIQAIAYhBgkCCEICUKCkCAECEIAghAAgBiEGCQIIQgJQoKQIAQIQgCCEACAGIQYJAghCAlCgpAgBAhCAIIQAIAYJAaJQYIQgpAghCAECEIAghAAgBgkBiEIIQgJQghCgCAEIAgBAGKQ4CIGIQghCAlCCEKAIAQgCAEAYhBikCAkCAlCpQxCnaiCUPLvCjCCECAIAQhCAABikBiEIIQgFHEQevBLfy7ACEKAIAQgCAEAiEFiEIIQgpAghCAECEIAghAAIAaJQWIQghCCkCCEIAQIQgCCEAAgBiEGIQghCAlCCEKAIAQgCBUo+SA+GI4AgH3qJwbhGo7GIpAYJAghCAlCgpAgBAhCAIIQNyNQq92brNVakzdXGwBAZJK/45O/66seh8QgQQhBSBAShAQhQBACEISqeb3N+sak2eoalAFAhSR/998avItBYpAghCBUcBB6KMgg9DMBRhACBCEAQSgmyTeEV9eaBmMAUEHJe4DBcCwGiUGCENUKQs8KQoKQIAQIQgCCkBgEAFRQrz8Ug8SgYAwFIUFIEBKEEIQAQQgQhEj3eUFiEABQhZNCYlC5YpAgJAgJQoIQghAgCAGCECmq1dsGYADAbbV6SwwiiBgkCAlChwtCY0FIEBKEAEEIQBDi3ZJrYQy+AIB36/YGYhCFxyBBSBAShAQhBCFAEAIEIVKyVmsZegEAd0neI4hBFB2DBCFBSBAShBCEAEEIEIRIwXA0NvACAHbVH4zEIAqNQcORICQICUKCEIIQIAgBghAza3f6hl0AwK7anZ4YRKExSBAShAQhQQhBCBCEAEGIFDSaHcMuAGBX9UZbDKLQGCQICUKCkCCEIAQIQoAgRAqSIY9hFwAQWxASg+KJQYKQICQICUIIQoAgBAhCCEIAgCAkBkUegwQhQUgQEoQQhABBCBCEEIQAAEFIDIo8BglCgpAgJAghCAGCECAIkYJmq2vYBQDsKnneoBhEkTFIEBKEBCFBCEEIEIQAQYgUdHsDwy4AYFftTk8MotAYJAhV16dO//wngpAgxJ5O2itAEAIQhNi35EO5YRcAsJvBcCwGUWgMGo7GglBFfXr5FytpBaGHBSFBSBACBCEAQQjPEQIAdrZWa4lBFB6DBCFBSBAShBCEAEEIEIRIyWA4MvQCAO6SXC0rBlF0DBKEBCFBSBBCEAIEIUAQwikhACAjyXsDMYgQYpAgJAgJQrMGoTVBSBACBCEAQYg7ksHK6lrTAAwAmL4nSAb5YhAhxCBBSBAShAQhBCFAEAIEIVKWfNgWhQBADBoMx2IQwcQgQUgQEoQEIQQhQBACBCEykHx4r9VdHwcAVVSrt8QggotBgpAgJAgJQghCgCAECEJkqN3pOy0EABU6FdTu9DwziCBjkCAkCBUdhG5GodCCUF0QQhACBCFAECLd5wr1+sPpQ6UNywAgPsnf8Z1uP+jnBYlBYpAgJAgJQoIQghAgCAGCEAUEosFwBACl1k8Mqu3WgL0UxCAxaPp6HQtCgpAgVEQQ+tCT/3PymW/9aPLFF5YmS4ufn5z93qOTU6f+2eTEC8uTT3zrTwUZQQgQhAAEIQAg0C83TL/gsN0GYhCBxyBBSBAShPINQh/72v+Y/KcfPD5547/9rclf/slfeYe/+MF73mGw/EuTc3MPTp588VvijCAECEIAghAAIAYhBolBh49BgpAgJAjlE4Q++wf/efLTP3rwrgi0VxDabm3pr05PD4k0ghAgCAEIQgCAGIQYJAYdOAYJQoKQIJRtEPrwU/9r8qMfPL5nCNpPENoehk68cEasEYQAQQhAEAIAxCDEIDFIEEIQCiEIHf+3Fye1V+/fVwzabxDa4rSQIAQIQgCCEAAgBiEGiUGCENUIQs+EG4SSGDS6+Mv7jkEHDUJ/cfY9k3OnHxRtBCFAEAIQhAAAMQgxSAwShBCEighCh4lBBwpCZ+8QhQQhQBACEIQAADEIMUgMEoQQhHIOQh9++n8f6Jq4Awehs3f75stfFG8EIUAQAhCEAAAxSAwSg8SgewWhdUFIEBKEUgpCr//oI4eKQfsKQmd3Nlj+pcknvvWnAo4gBAhCAIIQACAGiUFikBgkCCEIHT4I1fYVhD777T86dAy6ZxA6u7efLvwNAUcQAgQhAEEIABCDxCAxSAza3UgQEoQEoVSC0GGvirtnEDq7PydeOCPiCEKAIAQgCAEAYpAYJAaJQYIQglBWQWjW00G7BqGz+/ff594r4ghCgCAEIAgBAGKQGCQGiUGCEIJQVkHo1X//aPpB6OzB/cY3/p+QIwgBghCAIAQAiEFikBgkBglCCEJZBKHRxV9ONwidPZxvvvxFIUcQAgQhAEEIABCDxCAxRgwShBCE0g5CaVwX944gdPbwzp3+20KOIAQIQgCCEAAgBolBiEGCEIJQ2kHopbmvpReEzs7mpwt/XcgRhABBCEAQAgDEIDEIMUgQIuYg1C4kCJ1Z+lfpBKGz70mFkCMIAYIQgCAEAIhBYhBikCCEIBRiELoiCAlCgCAEIAgBAGIQYpAYJAghCMUbhK6kGISWBSFBCBCEAAQhAEAMEoMQgwQhBKGZg9D70wxCV1IMQsuCkCAECEIAghAAIAaJQYhBghCCUFhB6EqKQWhZEBKEAEEIQBACAMQgMQgxSBBCEAorCF1JMQgtC0KCECAIAQhCAIAYJAYhBglCCEJhBaErKQahZUFIEAIEIQBBCAAQg8QgxCBBiCCD0KC6QehKikFoWRAShABBCEAQAgDEIDEIMUgQQhAKKwhdSTEILQtCghAgCAEIQgCAGCQGIQYJQghCOQahz88cgw4UhJYFIUEIEIQABCEAQAwSgxCDBCEEobCC0JUUg9CyICQIAYIQgCAEAIhBYhBikCBEYUFoFF4QejqAIHQlxSC0LAgJQoAgBCAIAQBikBiEGCQIIQiFFYSupBiElgUhQQgQhAAEIQBADBKDEIMEIQShsILQlRSD0LIgJAgBghCAIAQAiEFiEGKQIIQgFFYQupJiEFoWhAQhQBACEIQAADFIDEIMEoQQhMIKQldSDELLgpAgBAhCAIIQACAGiUGIQYIQglBYQehKikFoWRAKwCv2ChCEAAQhAEAMQgwSg6KIQYJQdX3hh9cfE4RSDEJXUgxCy4JQIF63V4AgBCAIAQBiEGKQGBRFDBKEBKEwglBfENoKQsuzO/H8kpgjCAGCEIAgBABiEGIQYpAghCAUZBBaFoQEIUAQAhCEAAAxSAxCDBKEEITiDUKXBSFBCBCEAAQhAEAMEoMQgwQhBKF4g9BlQUgQAgQhAEEIABCDxCDEIEGIUgahoSB0gBgkCAlCgCAEIAgBAGKQGIQYJAghCMUYhC4LQoIQIAgBCEIAgBgkBiEGCUIIQvEGocuCkCAECEIAghAAIAaJQYhBghCC0L6C0AfKGIQuC0KCECAIAQhCAIAYJAYhBglCCELxBqHLgpAgBAhCAIIQACAGiUGIQYIQglC8QeiyICQIAYIQgCAEAIhBYhBikCCEIFTOILT4+ZljkCAkCAGCEIAgBABikBgkBiEGCUJkF4RuRSFBKMMgdFkQEoQAQQhAEAIAxCAxCDFIEEIQijcIXRaEBCFAEAIQhAAAMUgMQgwShBCE4g1ClwUhQQgQhAAEIQBADBKDEIMEIQShYoPQU2kFod+bOQYJQoIQIAgBCEIAIAYhBiEGCUIIQmUKQpcFIUEIEIQABCEAQAwSgxCDBCEEoXiD0GVBSBACBCEAQQgAEIPEIMQgQQhBKN4gdFkQEoQAQQhAEAIAxCAxCDFIEEIQijcIXRaEBCFAEAIQhAAAMUgMQgwShBCEBKE8gtAZQUgQAgQhAEEIAMQgxCAxSAwShBCE4g1CZwQhQQgQhAAEofCHgusbk8FwBEBF9BMDyqK3XX8vQw7gVogQgwQhBCFBKI0gdEYQEoQAQQhAEApWMrRotXuTWr09eXO1AQBQOWu15ub7oe40lIpBghCC0K5B6KQgtN8YJAgJQoAgBCAIBXYaKAlBhkAAAHc0W51DnxoSgwQhBKHKBqEzgpAgBAhCAIJQkJIP3Gu1lqEPAMAOVtea02v6xKD8DAQhQUgQKm8QOiMICUKAIAQgCAUbg5Ihh2EPAMDeOt2+GJRTDBKEBCFBqKRB6IwgJAgBghCAIBTs84LEIACA9E4KiUHpxCBBSBAShEoYhM4IQoIQIAgBCELBqjfahjsAAAdQq7fEoBxikCAkCAlCJQtCZwQhQQgQhAAEoWD1+kNDHQCAQ2i1e2JQxjFIEBKEBKESBaEzgpAgBAhCAIJQ0NZqLQMdAIBDWKs1xaCMY5AgJAjFH4RacQShM4KQIAQIQgCCUNCSD96GOQAAh9ftDcSgDGPQYCgICUKCUPBB6IwgJAgBghCAIBS8dqdvkAMAMNO1cV0xKMMYJAgJQoJQ4EHojCAkCAGCEIAgVAqNZscgBwBgBrVGWwzKMAYJQoKQIBRwEDojCAlCgCAEIAiVRr3RNsgBAJglCNVbYlCGMUgQEoTuGYSeE4QKCUJnBCFBCBCEAAQhQQgAoGLEoOxikCAkCAlCAQahM4KQIAQIQgCCkCAEAFDVE0JiUCYxSBAShAShwILQGUFIEAIEIQBByDOEAACq+gwhMSizGCQICUKCUEBB6IwgJAgBghCAIFRa3d7AIAcAYAbNVlcMyjAGCUKCkCAUSBC6JAgJQoAgBCAIlVrywdwgBwDg8JIv2IhB2cUgQUgQEoQCCEKXBCFBCBCEAAShKNTqniMEAHAYa7WmGJRxDBKEBKHqBaFmWEHokiAkCAGCEIAgFI3+YGSgAwBwCJ1uXwzKOAYNhiNBSBAShIoKQpcEocBds1eAIAQgCHFg9YZTQgAAB1Grt8SgHGKQIFRdJ//4+n2CUIFB6JIgVAb2ChCEAAQhDmy8vjFZXWsa7gAA7EPyvqnXH4lBOcQgQajaBKGCgtClbIPQqZcfF3MEIUAQAhCEipR8cBeFAADEoJBikCAkCAlCOQehS9kHobOnPi7mCEKAIAQgCIUQhWp118cBAOxkrSYG5R2DBCFBSBDKMQhdyiEILQlCghAgCAEIQkFpd/pOCwEAbNNsdafBQgzKNwZNg9BIEBKEBKHZgtCJmWNQKkFoSRAShABBCEAQCva5Qt3eYFJvODEEAFRTrd6aflGmP9jpVJAYlEcMEoQEIUEohyB0KYcgtCQICUKAIAQgCJXqOrm9PqgDkL1+YkBZ9Lbr72VIwbrv0ts1AIlBeccgQUgQCjcI9eIIQpdyCEJLgpAgBAhCAIIQAOz/5Ob09OZ2GwRstN14L+sUbLgTMSiYGCQICUKCUIZB6FIOQWhJEBKEAEEIQBACADFIDEIMEoMEIQShYoLQpRyC0JIgJAgBghCAIAQAYpAYhBgkBglCCELFBKFLOQShJUFIEAIEIQBBCADEIDEIMUgMEoQQhIoJQpdyCEJLgpAgBAhCAIIQAIhBYhBikBh0QENBSBAShNIJQpdyCEJLgpAgBAhCAIIQAIhBYhBikBgkCCEIFROELuUQhJYEIUEIEIQABCEAEIPEIMQgMUgQQhCKNwgtCUKCECAIAQhCACAGiUGIQWLQTEFoLAgJQoJQyEFoSRAShABBCEAQAgAxSAxCDBKDBCEEoXiD0JIgJAgBghCAIAQAYpAYhBgkBglCCELxBqElQUgQAgQhAEEIAMQgMQgxSAwShMgsCG0IQkUHoSVBSBACBCEAQQgAxCAxCDFIDBKEEITiDUJLgpAgBAhCAIIQAIhBYhBikBgkCCEIxRuElgQhQQgQhAAEIQAQg8QgxCAxSBBCEIo3CC0JQoIQIAgBCEIAIAaJQYhBYpAghCAUbxC6KAgJQoAgBCAIAYAYJAYhBolBghCCULxB6KIgJAgBghCAIAQAYpAYhBgkBglCCELxBqGLgpAgBAhCAIIQAIhBYhBikBgkCCEIxRuELgpCghAgCAEIQgAgBolBiEFikCCEIBRvELooCAlCgCAEIAgBgBgkBiEGiUGCEIJQvEHooiAkCAGCEIAgBABikBiEGCQGCUIEF4TWBaE9g9C/FIQEIUAQAhCEAEAMQgwSg8SgcGOQICQICUI5B6GLgpAgBAhCAIIQAIhBYhBikBgkCCEIxRuELgpCghAgCAEIQgAgBolBiEFikCCEIBRvELooCAlCgCAEIAgBgBgkBiEGiUGCEIJQmEHoyRSC0EVBSBACBCEAQQgAxCAxCDFIDBKEEITiDUIXBSFBCBCEAAQhABCDxCDEIDFIEEIQijcIXRSEBCFAEAIQhABADBKDEIPEIEEIQSjeIHRREBKEAEEIQBACADFIDEIMEoMEIQSheIPQxaKD0MfEHEEIEIQABCEAxCDEIDFIDBKDBCEEocyC0EVBSBACBCEAQQgAxCAxCDFIDBKEEITiDUIXBSFBCBCEAAQhABCDxCDEIDFIEEIQijcIXQwkCC0KQoIQIAgBCEIAiEGIQWKQGCQGCUIIQukHoYVAgtCiICQIAYIQgCAEgBiEGCQGiUFikCCEIBRvEFoUhAQhQBACEIQAEIMQg8QgMUgMEoQQhOINQouCUIaO2itAEAIQhABADBKDxCAxSAwqfQwShKrt159/a7AVhD4oCJUzCC0KQhk7Zq8AQQhAEAIAMUgMEoPEIDGo9DFIEKq2R0/9/A1BqMRBaHFn577/K0KOIAQIQgCCEABiEGKQGCQGiUGCEIJQ6YPQ4u5+OvfXhBxBCBCEAAQhAMQgxCAxSAwSgwQhBKF3BqFGuYLQoiAkCAGCEIAgBIAYhBgkBolBYpAghCAUbxBaFIQEIUAQAhCEABCDEIPEIDFIDBKEEITiDUKL+wxCpwUhQQgQhAAEIQDEIMQgMUgEEoMEIQSh8gWhRUFIEAIEIQBBCAAxCDFIDBKDxCBBiCKD0NcFoUyD0KIgJAgBghCAIASAGIQYJAaJQWKQIIQgFG8QWhSEBCFAEAIQhAAQgxCDxCAxSAwShBCE4g1Ci4KQIAQIQgCCEABiEGKQGCQGiUGCEJULQt3wgtBXMwpCi4KQIAQIQgCCEABiEGKQGCQGiUGCEIJQvEFoURAShABBCEAQAkAMQgwSg8QgMUgQQhCKNwgtCkKCECAIAQhCAIhBiEFikBgkBqWsLwgJQoJQCkHod9MJQouCkCAECEIAghAAYhBikBgkBolBGcQgQUgQEoQCCUIXBCFBCBCEAAQhAMQgxCAxSAwSgzKKQYKQICQIBRCELghCghAgCAEIQgCIQYhBYpAYJAZlGIMEIUFIECo4CF0QhAQhQBACEIQAEIMQg8QgMUgMyjgGCUKCkCBUYBC6IAgJQoAgBCAIASAGIQaJQWKQGJRDDBKEBCFBqKAgdEEQEoQAQQhAEKqs2AcQQGQDxQFl0duuv5chKRKDxKCyxCBBSBAShAoIQhcEIUEIEIQABKFKSQY/3d5gUqu3J2+uNgCAyNTqrUmr3ZsO48UgMSjUGCQICUKCkCCEIAQIQoAgRFbXLK1vTNqdvkEZAFRIq92dhgsxSAwKLQYJQoJQuYNQp3xB6IIgJAgBghCAIFQJydBirdYyGAOAClqrNafX+IlBYlBIMUgQEoQEoRyD0AVBSBACBCEAQagyMWh1rWkgBgAVlrwX2IpCYpAYFEIMSl6PgpAgJAjlEIQuCEKCECAIAQhClXlekBgEANyOQsmpDDFIDAogBglCgpAglEMQupBjEFoQhAQhQBACEIQKVW+0DcAAgNtq9ZYYJAYFEYMEIUFIEMo4CF3IMQgtCEKCECAIAQhCher1hwZfAMBdOt2+GCQGFR6DBCFBSBDKMAhdyDEILQhCghAgCAEIQoWr1Z0OAgDutlZrikFiUOExSBAShAShjILQhRyD0IIgJAgBghCAIFS4ZHhh4AUA7KbXH4lBYlChMUgQEoRyCULPhheEHsoyCF3IMQgtCEKCECAIAQhCQej2BoZdAMCuWu2eGCQGFRqDBCFBSBBKOQhdyDEILQhCghAgCAEIQsFoNDuGXQDArpKrZcUgMajIGCQICUKCUIpB6EKOQWhBEBKEAEEIQBAKSr3h+UEAwEGCkAgkBuUbgwQhQUgQSikIXcgxCC0IQoIQIAgBCEKCEABQ4iAkAolB+ccgQUgQOnwQGgtCRQShBUFIEAIEIQBBSBACAEochEQgMaiYGCQICUKCUImC0MJ+g9D9Qo4gBAhCAIKQZwgBAOEFIRFIDCouBglCgpAgVJIgtCAICUKAIAQgCAWt2xsYdgEAu2q1u0KQGFRoDOoPhoKQICQIhR6EFgQhQQgQhAAEoeAlww3DLgBgN73+UAwSgwqNQYKQICQIpRGEPpddEFoQhAQhQBACEIRKI7kKxsALAHi3tVpTDBKDCo9B0yA0FIQEIUEoyCC0IAgJQoAgBCAIlUryzV9DLwDg3TrdvhgkBhUegwQhQUgQCjQILQhCghAgCAEIQqVUbzglBADcUau3xCAxKIgYJAgJQoJQgEFoQRAShABBCEAQKq3ReH2yutY0AAMApu8JksG8GCQGhRCDBCFBSBAKLAgtCEKCECAIAQhCpZcMP0QhABCDkutkxSAxKJQYJAgJQoJQQEFoQRAShABBCEAQiioK1equjwOAKlqriUFiUHgxKDEQhCrrU6d//hNBKJAgdD7FIPR9QShFJ+0VIAgBCEIc2nh9Y9Lu9A3GAKBCmq3udOAvBolBocUgQajaPr38i5W0gtDDgtBMMSjNIPR/5+4TcgQhQBACEIRCe65QtzdwYggAIlWrtyatdrfyzwsSg8KOQYKQICQIFRyEzqcfhBJCjiAECEIAglDAYh90ADkNFAeURW+7/l6GFKy7k97eqh6AxKDyxCBBSBAShAoMQucFIUEIEIQABCEADnod5fRKyu02CNhou/Fe1inYcCejexGBxKDyxCBBSBAShNIIQr87cwwShAQhQBACEIQAEIPEIMQgMUgMyiwGCUKCkCBUQBA6LwgJQoAgBCAIASAGiUFikBgkBolBOcagm0FoJAgJQoKQIIQgBAhCgCAEgBiEGCQGiUFiUKwxSBAShAShnIPQeUFIEAIEIQBBCAAxSAwSY8QgMUgMyjkGCUKCUAhB6GYUCi0I1dMPQucFIUEIEIQABCEAxCAxSIwRg8QgMaiAGCQICUKCUE5B6LwgJAgBghCAIASAGCQGiTFikBgkBhUUgwQhQUgQyiEInReEBCFAEAIQhAAQg8QgMUYMEoPEoAJjkCAkCAlCGQeh84KQIAQIQgCCEABikBgkxohBYpAYVHAMEoQEIUEowyB0XhAShABBCEAQAkAMEoPEGDFIDBKDAohBgpAgJAhlFITOC0KCECAIAQhCAIhBYpAYIwaJQWJQIDFIEBKEBKEMgtB5QUgQAgQhAEEIADFIDBJjxCAxSAwKKAYJQoJQ6YPQM4EFofOCkCAECEIAghAAYpAYJMaIQWKQGBRYDBKEBCFBKMUgdD6QIDQvCAlCgCAEIAgBiEGIQWKQGCQGiUGCEIJQ+kHofCBBaF4QEoQAQQhAEAIQgxCDxCAxSAwSgwQhBKFDBqFa+EFoXhAShABBCEAQAhCDEIPEIDFIDBKDBCEEoYCD0JHUYpAgJAgBghCAIAQgBiEGiUFikBgkBglCCEKpB6HPzRyDZgpC84KQIAQIQgCCEIAYhBgkBolBYpAYJAghCAUchI7MFoTmBSFBCBCEAAQhADEIMUgMEoPEIDFIEEIQCjgIHZktCM0LQoIQIAgBCEIAYhBikBgkBolBYpAghCAUcBA6MlsQmheEBCFAEAIQhADEIMQgMUgMEoPEIEEIQSjgIHRktiA0LwgJQoAgBCAIAYhBiEFikBgkBolBghCCUMBB6MhsQWheEBKEAEEIQBACEIMQg8QgMUgMEoMEISofhNoBB6EjswWheUFIEAIEIQBBCEAMQgwSg8QgMUgMEoQQhIoJQvOfmzkG3TMIzQtCghAgCAEIQgBiEGKQGCQGiUFikCCEIBRwEDoyWxCaF4QEIUAQAhCEAMQgxCAxSAwSg8QgQQhBKPcg9P59B6EjswWheUFIEAIEIQBBCEAMQgyfSchzAAAgAElEQVQSg8QgMUgMEoQQhAIOQkdmC0LzgpAgBAhCAIIQgBiEGCQGiUFikBgkCCEIBRyEjswWhOYFIUEIEIQABCEAMQgxSAwSg8QgMUgQQhAKOAgdmS0IzQtCghAgCAEIQgBiEGKQGCQGiUFikCBEFEFoEGkQOjJbEJoXhAQhQBACEIQAxCDEIDFIDBKDxCBBCEEo4CB0ZLYgNC8ICUKAIAQgCAGIQYhBYpAYJAaJQYIQglDAQWi2GPSX5wQhQQgQhAAEIQAxCDFIDBKDxCAxSBBCEDpcEHq6BEHonCAkCAGCEIAgBCAGIQaJQWKQGCQGCUKUJgiNBKFDxiBBSBACBCEAQQhADEIMEoPEIDFIDBKEEIRiDELnBCFBCBCEAAQhADEIMUgMEoPEIDFIEEIQijcInROEBCFAEAIQhADEIMQgMUgMEoPEIEEIQSjeIHQu2yB0QxAShABBCEAQAhCDxCAxSAwSg8QgMWi7niAkCAlCUQWhG4KQIAQIQgCCEIAYJAaJQWKQGCQGiUHvjkGCkCAkCOUchM5lF4RuCEJZeMVeAYIQgCAEIAYJLmIQYpAYJAaVPgYJQtX2hR9ef0wQyjEIncsuCN0QhLLyur0CBCEAQQhADEIMQgwSg8Sg0scgQUgQCicI9eMOQueyC0I3dnDi+TkxRxACBCEAQQhADBKDxCAxSAwSg8QgQQhBKLcgdC67IHRDEBKEAEEIQBACEIPEIDFIDBKDxCAx6F4xSBAShAShjIPQueyC0A1BSBACBCEAQQhADBKDxCAxSAwSg8Sg/cQgQUgQyjYIDasdhM5lF4RuCEKCECAIAQhCAGKQGCQGiUFikBgkBu03BglCgpAglFEQOpddELohCAlCgCAEIAgBiEFikBgkBolBYpAYdJAYJAgJQoJQBkHoXHZB6IYgJAgBghCAIAQgBolBYpAYJAaJQWLQQWOQICQICUJpBKHPzhyD9hOEbhwkCH1bEBKEAEEIQBACEIPEIMQgMUgMEoMEISIKQh8IJQidyy4I3RCEBCFAEAIQhADEIDFIDBKDxCAxSAw6bAzq9QUhQUgQSiUIncsuCN0QhAQhQBACEIQAxCAxSAwSg8QgMUgMmiUGCUKCkCAUdhC6IQgJQoAgBCAIAYhBYpAYJAaJQWKQGDRrDBKEBCFBKNwgdEMQEoQAQQhAEAIQg8QgMUgMEoPEIDEojRgkCAlCtwffglBQQejGzEHotJgjCAGCEIAgBCAGiUGIQWKQGCQGCUIIQqEGoRuCkCAECEIAghCAGCQGiUFikBgkBolBacYgQUgQEoTCCkI3BCFBCBCEAASh+E0HQZEPciCYgeKAsuht19/LkIJ1d9K7lwGp6ZdKrz8QgwKJQYKQIFT5IPRUOEHohiAkCAGCEIAgFOkJhfWN6QCn3mhP3lxtAABUzlqtNWm1e1tRQgwqIAYJQoKQIBRGEHpbEBKEAEEIQBCKMwS1O/3J6lrTIAgA4JZmqzMNHWJQvjFIEBKEBKHig9DbgpAgBAhCAIJQnNfC1epOBAEA7HxiqHn7OjkxKJ8YJAgJQoJQsUHobUFIEAIEIQBBKM4Y5FQQAMDekvdL3f5ADMopBglCgpAgVFwQelsQEoQAQQhAEIrzmjgxCAAgxSgkBqUSgwQhQUgQKiYIvTsGvf2qICQIAYIQgCAUhXrDNXEAAAe7Pq4lBuUQgwQhQUgQyj8I7RSDBCFBCBCEAAShCCRDCEMdAICDa3V6YlDGMejWM5sEIUEo/CB0Mo4gtFsMEoQEIUAQAhCEIlCrOx0EAHCoq+NqTTEo4xgkCAlCglB+QWivGCQICUKAIAQgCJXccDQ2zAEAmEG72xeDMoxBgpAgJAjlE4TuFYMEIUEIEIQABKGS6/YGBjkAADNotDpiUIYxSBAShASh7IPQfmKQICQIAYIQgCBUco1mxyAHAGAGtXpLDMowBglCgpAglG0QelsQEoQAQQhAEKqGesPzgwAA8gtCYtBBY5AgJAgJQtkFoYPEIEFIEAIEIQBBSBACAKg8MSi7GCQICUKCUDZB6KAxSBAShABBCEAQEoQAACptrdYSgzKMQYKQIFSNINTKNQgdJgYJQoIQIAgBCEKeIQQA4Mo4MSizGCQICUKCULpB6LAxSBAShABBCEAQKrl2p2+QAwAwg+QLNmJQdjFIEBKEBKE0gtBnZo5BgpAgBAhCAIJQyQ1HY4McAIAZJF+wEYOyi0GCkCAkCKUThGaNQYKQIAQIQgCCUASSe+8NcwAADm51rSkGZRyDBCFBaF9B6DlB6MBB6FVBSBACBCEAQahykg/lBjoAAAfXbHXFoIxjkCAkCAlCGQShVwUhQQgQhAAEocqqN9qGOgAAB5CcshaDso9BgpAgJAilHIReFYQEIUAQAhCEKm00Xp9eeWK4AwCwv6viur2BGJRDDJoGoYEgJAgJQqkEoVcDCUJzgpAgBAhCAIJQoYajsSgEALAP7U5fDMopBglCgpAglFIQejWQIDQnCAlCgCAEIAgFE4WS608MegAAnAwKIQYl+oKQICQIxRGE5gQhQQgQhAAEoaCM1zcmrXbP0AcAYJt6ozMNHGJQvjFIEBKEBKFIgtCcICQIAYIQgCAU9HOFkutQavW2IRAAUNkTQY1mZ9LtvTsEiUF5xSBBSBCqZhBqxhWE5gQhQQgQhAAEoVKdGhoMR1Bp/eFoh2Egoept19/LkIJ1d9K7lwGp6Uets1/du919GkgMKiIGCUKCkCBU8iA0JwhlbGSvAEEIQBACSDOKTsPodhsEbLTdeC/rFGy4k9G9jLllsJvhflUg5O/HgaOzGJRnDBKEqu3kH1+/TxAqcRCaE4TyYK8AQQhAEAIQg8QgMUgMEoPEIDGo9DFIEEIQKmkQmtvbqRf/kZgjCAGCEIAgBIhBiEFikBgkBolBYpAghCBU2iA0d29nX/4HYo4gBAhCAIIQIAYhBolBYpAYJAaJQYIQglApg9CcICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEIBRvEJoThAQhQBACEIQAMQgxSAwSg8QgMUgMEoSILgj1BKFDxCBBSBACBCEAQQgQgxCDxCAxSAwSg8QgQQhBqGxBaE4QEoQAQQhAEALEIMQgMUgMEoPEIDFIEEIQijcIzQlCghAgCAEIQoAYhBgkBolBYpAYJAYJQghC8QahOUFIEAIEIQBBCBCDEIPEIDFIDBKDxKDUgtBQEBKEBKHQgtCcICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEIBRvEJoThAQhQBACEIQAMQgxSAwSg8QgMUgMEoQQhOINQinEoBunBSFBCBCEAAQhQAxCDBKDxCAxSAwSgwQhBKF0g9BcSkEopRgkCAlCgCAEIAgBYhBikBgkBolBYpAYJAghCIUYhH58JLUYJAgJQoAgBCAIAWIQYpAYJAaJQWKQGCQIIQiFFoR+nEIQOi0ICUKAIAQgCAFiEGKQGCQGiUFikBgkCCEIhRmEfpxCEDotCAlCgCAEIAgBYhBikBgkBolBYpAYJAhxqCC0IQhlHYR+nEIQOi0ICUKAIAQgCAFiEGKQGCQGiUFikBgkCCEI5RCE/sXMMehQQei0ICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEIBRmEPpxCkHotCAkCAGCEIAgBIhBiEFikBj0/9m7syC7qzvB861mOmK27q4ZPehtoueBmJkXoqNdFUE4YqYWasozqqnqmqroQSC3oWwWG6mqELIN2ELYBhsDlrVLCBCIrTBFagW33RZbTZdtZNksUi439+XmzT2TRdiKqX74z/2nlFJKyuWu//s///t5+ETYSIjMezNv3nO++p0jBolBYpAghCCUziD0Sg2C0B5BSBACBCEAQQgQgxCDxCAxSAwSg8QgQQhBKLtBaI8gJAgBghCAIASIQYhBYpAYJAaJQWKQIIQglN4g9EqVQWiPICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEIJTeIPRKlUFojyAkCAGCEIAgBIhBiEFikBgkBolBYpAghCCU3iD0SpVBaI8gJAgBghCAIASIQYhBYpAYJAaJQWKQIIQglN4g9EqVQWiPICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEIJTeIPRKlUFojyAkCAGCEIAgBIhBiEFikBgkBolBYpAghCCU3iD0SpVBaI8gJAgBghCAIASIQYhBYpAYJAaJQWKQIETiQehjQajUIPRKlUFojyAkCAGCEIAgBIhBiEFikBgkBolBYpAghCCU3iD0SpVBaI8gJAgBghCAIASIQYhBYpAYJAaJQWKQIIQglN4g9EqVQWiPICQIAYIQgCAEiEGIQWKQGCQGiUFikCCEINSYILSphCBUZQz6x2OCkCAECEIAghAgBiEGiUFikBgkBolBghCCUHaD0DFBSBACBCEAQQgQgxCDxCAxSAwSg8QgQQhBKLtB6JggJAgBghCAIASIQYhBYpAYJAaJQWKQIIQglN0gdEwQEoQAQQhAEALEIMQgMUgMEoPEIDFIEEIQym4QOiYICUKAIAQgCAFiEGKQGCQGiUFikBgkCCEIZTcIHROEBCFAEAIQhAAxCDFIDBKDxCAxSAwShBCEshuEjglCghAgCAEIQoAYhBgkBolBYpAYJAYlbFIQEoQEoeSC0DFBSBACBCEAQQgQgxCDxCAxSAwSg8SgBsQgQQhBKKEgdCzpIPSnYo4gBAhCAIIQiEFikBiEGCQGiUFikBgkCCEIJRaEjglCghAgCAEIQoAYhBgkBolBYpAYJAY1MAYJQghCtQhCX6o6BglCghAgCAEIQoAYJAaJQWKQGCQGiUFiUN1ikCCEIFTHIHRMEMqIf+W1AgQhAEEIEIMQg8QgMUgMEoPEoKBjkCDEn3zvk5m5IPQHglDtgtAxQShDfs9rBQhCAIIQIAYhBolBYpAYJAaJQUHHIEGI63f8OicI1TgIHWt8EHpr5/8s5AhCgCAEIAiBGIQYhBgkBolBYpAYJAghCNUlCB1LRxA6ufN/EHIEIUAQAhCEQAxCDEIMEoPEIDFIDBKEEIQuDUIj1QehY4KQIAQIQgCCECAGIQaJQWKQGCQGiUEpjEGCEIJQjYLQMUFIEAIEIQBBCBCDEIPEIDFIDBKDxKCUxiBBCEEoo0FohyAkCAGCEIAgBGIQYhBikBgkBolBYpAghCCU3SC0WxAShABBCEAQAjEIMQgxSAwSg8QgMWi+KUFIEKpREHpAEEpFENotCAlCgCAEIAiBGIQYhBgkBolBYpAYdFkMEoQQhDIUhHYLQoIQIAgBCEIgBiEGIQaJQWKQGCQGLRCDBCEEoYwEod2CkCAECEIAghCIQYhBiEFikBgkBolBi8SgyalpQUgQCiwITaYvCD3W4CC0WxAShABBCEAQAjEIMQgxSAwSg8QgMWiJGCQIIQgFHoR2C0KCECAIAQhCIAYhBiEGiUFikBgkBi0TgwQhBKGAg9BuQUgQAgQhAEEIxCDEIMQgMUgMEoPEoBJikCCEIBRoENotCAlCgCAEIAiBGIQYhBgkBolBYpAYVGIMEoQQhAIMQrsFIUEIEIQABCEQgxCDEIPEIDFIDBKDyohBghCCUGBBaLcgJAgBghCAIARiEGIQYpAYJAaJQWJQmTFIEEIQCigI7RaEBCFAEAIQhEAMQgxCDBKDxCAxSAyqIAYJQghCgQSh3YKQIAQIQgCCEIhBiEGIQWKQGCQGiUEVxiBBCEEogCC0WxAShABBCEAQAjGIpohB8UZ8vKk3Nj51iYnJ6dlN6LRFl/hjWujjjf9ZIz9eMUgMEoPEIDFIEEIQCi4I7RaEBCFAEAIQhEAMIvMxKN7sHBmdiAaHRpaUHx6NxiemZzftGxmC4kA1XBhb9uONf0/8e8UgMUgMEoPEoMbHoNiUICQICULpDEK7BSFBCBCEAAQhEIPIdAyKN5gLI+PLhpWFwlC8CZh0CIo3rksJQQuFofjfFYPEIDFIDBKDGheDBCHCD0IT2QxCuwUhQQgQhAAEIRCDyHQMijc6h/KjZceV+cbGJxOdCqrmY43Vc1pIDBKDxCAxSAwShBCEggtCuwUhQQgQhAAEIRCDyHwMqjauzBkdmwgiBtUzColBYpAYJAaJQYIQglBwQWi3ICQIAYIQgCAEYhCZPyau2smgJKNQLWPQnHizVwwSg8QgMUgMSjYGCUIIQikKQrsFIUEIEIQABCEQg8h0DIpVcmdQo6JQPWLQ3B1IYpAYJAaJQWJQsjFIEEIQSkkQOioICUKAIAQgCIEYROZjUC2Piqt3FKpXDJozPjEtBolBYpAYJAYlGIMEIQShFASho4KQIAQIQgCCEIhBZD4G1XM6qNZRqN4xqNopITFIDBKDxCAxSBBCEAouCB0VhAQhQBACEIRADKIpYlC8EV/vyFKLKJREDJoTb5KLQWKQGCQGiUHJxCBBiMSC0LfSF4T+t5oFoS9WHYMEIUEIEIQABCEQg8hwDIrFm3pJhZZKo1CSMSg2Nj4lBolBYpAYJAYlFIMEIQShBgWho4KQIAQIQgCCEIhBNE0MisXxI8nYUm4USjoGlfvxiUFikBgkBolBghCCUHBB6KggJAgBghCAIARiEE0VgxoVhEqNLo2IQbH4TiUxSAwSg8QgMSiZGDQbhKYFIUFIEEosCB0VhAQhQBACEIRADKLpYlAjg9ByUahRMajUICQGiUFikBgkBglCpCEIfSQIlROEjiYUhHYJQoIQIAgBCEIgBpGqGNToILRYFGpkDColCIlBYpAYJAaJQYIQglBwQehoQkFolyAkCAGCEIAgBGIQqYtBsfGJxsaXy6NQo2NQLI5kYpAYJAaJQWJQMjFIEEIQSiAIHU0oCO0ShAQhQBACEIRADCKVMSgWbxY3OsDMRaE0xKBYvAEqBolBYpAYJAYlE4MEIQShOgehowkFoV2CkCAECEIAghCIQaQ2Bs3JD4+mIsSkRRwvxCAxSAwSg8Sg6QSD0IwgJAgJQvUIQkcTCkK7BCFBCBCEAAQhEINIfQxKwz1CabLQnUZikBgkBolBYpAghCAUXBA6mlAQ2iUICUKAIAQgCIEYRBAxaDZ4fPhRNJQ3JRSLN+jFIDFIDBKDxCBBCEEo6CB0NKEgtEsQEoQAQQhAEAIxiGBi0Jx4E7DZY1A8KSUGiUFikBgkBglCCEJBB6GjCQWhXYKQIAQIQgCCEIhBBBeD5sTHpTVrDBoZnRCDxCAxSAwSgwQhBKGwg9DRhILQLkFIEAIEIQBBCMQggo1BzRyFhgtjsxFDDBKDxCAxSAwShBCEgg1CRxMKQrsEoQb4M68VIAgBCEIgBolBYpAoJAaJQWKQGCQGBR2DBCE+u+fXJwWhQILQLkGoQb7htQIEIQBBCMQgMUgMEoXEIDFIDBKDxKCgY5AgxBf3/+ZArYLQ7wtC9QtCu8oztPOfCzmCECAIAQhCIAaJQWmPQc0QhcQgMUgMEoPEoGlBCEFIECotCO2qjJAjCAGCEIAgBGKQGBRADMpyFEpDDHr+hR9Ef/wnfxH9T//Lv15Q/Gtrbrg5euR726Ijx16N8sOFTMSgoXwhOnL01eiRR7dF1xc/v9/9/c8s+hjM+dRvf7r4e2+K7rv/gei54uPW1pHLTAw6/vpb0cOPbo1uuW1ddP2NNy37WMx9bdxy67rZf+/4a29mJga1tndEzz7/YrRp8wPRmhs/t+TXxhduuyP6SfFzF4OyEYMEIQShlAehXYKQIAQIQgCCEIhBZD4GZTEKNToGnfjFL5cMQUuJA9GefftTFYdKiUFtHZ3R3sf2V/x5LySOBXEgevvEyeBi0OGjr0YbNt4d/Zvf/nTNHo9bbr0jeu75F4tf4/mgYlAcgeIAVOnXRhyGBgbzYlDgMUgQQhBKcRDaJQgJQoAgBCAIgRhE08SgLEWhRseg9o7O6FO/U5sIsGHjPdHrb7yV6hj02utvRbfetr5m0WOpiZl4cijNMWgwPzw70VPLCLSQ+M+/b/MDUVt7R6pjUDwJFE8B1er5F4PCjkGCEIJQSoPQLkFIEAIEIQBBCMQgmi4GZSEKpeGYuHjCp9YBIP4z46mjNMWgOARdX4fPtZSpobSEoaRD0ILR8K67UxeGDh15paRjAsv18CNbxaCAY5AghCCUwiC0SxAShABBCEAQAjGIpo1BIUehNMSgeJqnnpv/m+9/MLGj5BaLQfH9QPHkUtLhY6GJkThKNToG7XnsyYaEoMsnhuIg1egQ9PO3T9ZsImixz3NgcEgMCjQGCUIIQksFoUJpQWhvDYPQLkFIEAIEIQBBCMQgmj4GhRiF0hCDYkmEkvg4uiPHXm1IDIoncz7V4PhxufiOoaH8cOIxqK0jF11/w02peiziSBZHmUbEoDhIJfE5Pvvci2JQoDFIECItQehcFGryILRLEBKEAEEIQBACMQgxKMAolJYYVK/j4pa6X6ge00ILTgUV/ztJ3BNUTQh5+8TJxGJQHMb+TcrC2Hx79j6RWAiKj6uLH/+kPreHH/m+GBRoDBKEEIRSEoSOCEKCECAIAQhCIAYhBgUYhdIUg5IOQnMhpJZ3Cy0Ug94u/vn1uA+mHup9t1B8V9CGjXcH8Vjccusdxe+RfF1j0OEjryQexrIahJohBglCCEK1CEK3Vx2DBKFUu9lrBQhCAIIQiEGIQaJQADGoEUFo7gi551/4QV1i0N59+4OIH/Pdetu6uhwh9/MTJxOdhKmFOOQdf+3NusSg+zY/0JDPKYtBqFlikCCEINTgIHREEEqxgaLf8zoBghCAIARiEGJQKkxMTqcuCI2MTqQqBiV1h9CiEyG3r6/4CLmFjoi7vgFxq5Yh5LXX36pZDNrz2JPBPhazEeXRrTULQfEdRY0MY1m7Q6iZYpAgxDcOnl01G4UEoeSD0BFBKMW2Ff2W1wgQhAAEIRCDEIPEoGXEk0tpiUGxI8debejGfyXTQgtNBcV/TsgBZM599z9Q1bRQfC/R9TfclInHIo441UwLxcfPxWGp0Z/HwOCQGBRoDBKEmHPvD85e9+dbP8kLQgkFoSOCkKkgQBACEIRADEIMCjwGXZgUujwKNSgGNfLYuIUmZOIw1N7RWVIMaiv+vjgEhXJXUFmR7Lc/PRuG4rhTagg6cvTV2aPnsvZYxK6/8XPRc8+/WPL9QvFEUByCkr4rKOvHxTVjDBKEuNzt+39zQBCqcxA6IgiZCgIEIQBBCMQgxKCMxKArolCDY1AsjjBpmrCJI08cqTbf/2D0yPe2XXBf8f/Hx8JlMQItFYfiiZ8NG++OHnl06yXiABTaHUG1mBqKA1EcfObbcNfds/88DRHo4sf655mZDmrWGCQIsZCv/93Za/6f7Z/kgglC9wcUhI4IQqaCAEEIQBACMQgxKGMxaP6dQo2OQXNO/OKXTRVaoJ7W3PA5MSgDMWhCEGIJ657+9dbPPHTmrCBUoyB0RBAyFQQIQgCCEIhBiEEZjUHLR6GPEpcfLkR79u1vuqkTqJUv3LYueva5Fx0Tl5EYJAix7LTQS7+5Zu2uT04KQlUGoSOCkKkgQBACEIRADEIMyngMWjwKfZQK8dTQ62+8NevIsVdnj2275fb1TXFMW3wcW3wsW3w3z2uvv3WF+NfiY9yaYaoqDoT3bX5g9h6f46+9eYX4n8fHtsVHtmX9sYiPpLvzrrtn7wb6yWtvXNDa1p6ZCCQGXYxBghCl2vDsr9d95qGPzzZ3EBquLAgdEYRMBQGCEIAgBGIQYlCTxKAro9BHqRdPEj3/wg8yF0Piz+e54uc188GHZYkDUXzPT9bCRxyB2to7oumZD0oW//44DqXpLp9aHQF36PAr0dT0B5kLP2LQ4jFIEKIcm1/+zaobd505KQiVEYSOCEKmggBBCEAQAjEIMajJYtClUeijoMRTQ1mYCNr72JNlh6CFwlAWIlk86VNuCLrc4FA+uuXWOzIRxi6GIDGo2WKQIEQlvvz8r9f88SMfzwhCywShI4KQqSBAEAIQhEAMQgxq0hgUchSKj5YL9d6h+ON++8TJqmPQnKH88OxRcqHGjz17n6gqBF3u8JFXgp0W+sJtd0QDg3kxqIljkCBEpe57+derPr/vk8OC0CJB6IggZCoIEIQABCEQgxCDmjwGhRyF4mPkNmy8J6gN//vuf6BmIehy8d1DnwoohMRh7Odvn6xpDJo/LRTa/UK79zwxLwSJQc0agwQhqrXx+U/W/PEjH80IQtXFIEHIVBAgCAEIQiAGiUFikCiUQvHdQp/6nU+n/oi4ONjUKwbNaevIBTE5teGuu+sSgi4X3y2U+nukfu8z0c/ePikGiUGCEDV12xNnDghClccgQchUECAIAQhCIAaJQWKQKOQIufLvx7nhptlQU+8YNF88iZTWI+LiI92SiEFzjr/2ZmqPkLvyiDgxqNljkCBELX31hU+u+7MtH+WbNggdSVEQ2vlPTQUBCEIAghBiEGKQGJQ+o2OTQUah2CPf25aqqaC9jz2ZaAia77XX34p+9/c/k54wduNNUVt7R6IxaP4RcvFUUprC2KHDr1wWgsQgMUgQoj5uffzjA3/0nQ/PNlUQOpKiILSzKYPQe6aCAEEIQBBCDEIMCsL0zIdNG4PmxJuvoUah9o7OaM0NNzd0w//W29YlPhW0kKH8cPTIo1sberdQHKUOH3m1ISFooWmhRk+Sbdr8wAJTQWKQGCQIUV/3vPjJNf9u60e5xgSh8eYNQjubMgh9w/ccIAgBCEKIQYhBwcgPjzZ9EBrKj84GhVCjUOz1N95KPAzFx8PFkzmNDkEL3S20YePdiYeg557/wWxgTUMMmu+5519MfHrqzrvujlrbOhYIQWKQGCQIkZwvPvnx1j/69gdnBaEEgtDOpgtC8VTQv/Z9BghCAIIQYhBikKPiAjQ2Phl0EJofhjZsvKeuR8PFseXtEydTF4IWmxiqZwyJj4a7GILSF4Pmi+8zuuXWO+p6NFw8EbR4CBKDxCBBiORtemoMuVMAACAASURBVOmTVTfs+OikIFTHILSz6YKQqSBAEAIQhBCDxCAxKDzDhTExaN6UUBaCUGymaGi4ED33wg+iW29fH33qdz5d9fRLHIHiPy+OLGkPQQuJA9Z99z9QkyPU4gi0Z++TUVt7bl4ISncMmi++22jP3idqEod+9/c+MxuBFr4jSAwSg5YxKQiRnL85cGbd/x5PC2UkCP2vaQlCO5sqCJkKAgQhAEEIMUgMEoPCFG+SpyHExFFqZHTCXUI1jEELaevojI4cfTV65NFtsxNE199w8yJumg0n8WRN/PvTcDdQLU3HX/f54ej4629FDxc/x1j8OV/hxnNuuXXd7O+Jp4COv/bWZQEovBi0kJ+/fTJ69vkXZz/P+Ki3NTd+blFx/Hn4ka3RT157c5G7gcQgMaj0GCQIkbSvv3Rm1Wd3ffSGIFSjILSzqYKQqSBAEAIQhBCDxCAxyHFx1cagOGLEH8/o2IRj4+oUg2Y+KNWHmTZdqplyfRC0qXJMV0IMEoMWjkGCEI2y4dmP16z+7syMIFRFENrZNEHIVBAgCAEIQohBYpAYFL6x8anUxKDYB0UjDY5ChZFxMUgMEoPEIDEooRgkCNHQaaEfnFl1854PDwtCFQShnU0ThEwFAYIQgCCEGCQGiUGCUD1i0AcpiELDhXExSAwSg8QgMSihGCQIkYppoWc+XvNvH53JC0K1i0EZCEKmggBBCEAQQgwSg8QgQajeMehCFGrQnUIhBiExSAwSg8SgUGOQIESafOGxDw8IQrWJQYEHIVNBgCAEIAghBolBYpAglFQM+uDDcxoRhUI7Mk4MEoPEIDEo5BgkCJE2G5/7+Lo/vWRaKIQgdFsyQWhn5oOQqSBAEAIQhEAMEoOyK96IS2sMalQUGhufFIPEIDFIDBKDEopBghBpddvjH279wwenz9YkCG3OQBDamfkgZCoIEIQABCEQg8SgbIs3zdMcgxoRheINWzFIDBKDxCAxKJkYJAiRZl95/uNr/mLLdK7pg9DOTAchU0GAIAQgCIEYJAY1jzjUpDkGJRmFhvKjYpAYJAaJQWJQgjFIECIEX3ryw81/+ODU2aYMQjszHYRMBQGCEIAgBGKQGOTYuLTFoLkQUu8oFMJxcWKQGCQGiUFZikGCEKG4928/WnX91umTTRWEdmY2CJkKAgQhAEEIxCAxqHnlh0dTH4PqHYXi6aA4KIhBYpAYJAaJQcnFIEGI0Kx/6sN1f/jA5NnMB6GdmQ1CpoIAQQhAEAIxSAxqbvGmbggxqJ5RKN6UFIPEIDFIDBKDko1BghAhuueFj1Z9btfM4cwGoZ2ZDEJvFf0rX7+AIAQgCIEYJAZR46Pj6hmD6hGF4j9LDBKDxCAxSAxKPgYJQoTsr5/+YM3/+e3JmUwFoZ2ZC0IfFt3p6xUQhAAEIRCDxCDqEIXm4ko9Y1Ato5AYJAaJQWKQGNS4GCQIEf600IerPrdr+nAmgtDO2gahP30oZyoIQBACEIQQgxCD0n58XKV3Co2NT13yZ9UzBs2JNxPj+38quTPIMXFikBgkBolBjY1BghBZseHAB9f9yXcn88EGocO1D0J3PrLTVBCAIAQgCCEGIQalXRwj4rhTamgZHZuY3aBPOgZdCCfF/3Y86VPKxxv/ntGxydl/RwwSg8QgMUgMamwMEoTImr/cM30guCB0OFNByFQQIAgBCEIgBolBVDMxFMehOLgURsYvGBufvDBhc0VQSjAGXR6G4k3Z+GMbLoxfIv5n8a+lOQKJQWKQGCQGNVsMEoTIojsPfHDdnz86mQsiCB2uZxDaYSoIQBACEIQQgxCDMj1d1KAYlBVikBgkBolBzRSDJianBCEy65a901uv++b42dQGocOZCUKmggBBCEAQAjFIDEIMEoPEIDFIDBKD0hyDBCGybuMzH1zzfz86kUtdEDqciSBkKggQhAAEIRCDxCDEIDFIDBKDxCAxKIQYJAjRLG7fN735um+OnU1FEDqciSBkKggQhAAEIRCDxCDEIDFIDBKDxCAxKJQYJAjRTL763Myqf7dl4mRDg9Dh4IOQqSBAEAIQhEAMEoMQg8QgMUgMEoPEoNBikCBEM/rSE9Pr/o8Hx2YSD0KHgw9CpoIAQQhAEAIxSAxCDBKDxCAxSAwSg0KMQYIQzeorz82s+uyOycOJBaHDCQehHTUNQqaCAEEIQBACMUgMQgwSg8QgMUgMEoNCjkGxSUGIJrb+yek1n3lgdKauQehwwkFoR02DkKkgQBACEIRADBKDEIPEIDFIDBKDxKDQY5AgBNE/+cqz06tu2jl5oC5B6HDCQWhHzYKQqSBAEPIgAIIQiEFikBgjBolBYpAYJAaJQVmJQYIQXPTXT01f9399ZyxfsyB0OOEgtKNmQchUEIAgBAhCIAaJQWKMGCQGiUFikBgkBmUpBglCcKWbdk4cqDoIHU44CO2oSRAyFQQgCAGCEIhBYpAYJAaJQWKQGCQGiUFZjEGCECzszqenr/mzh8dyFQWhwwkHoR01CUJHin7Lcw8gCAGCEIhBYhBikBgkBolBYpAYlMEYJAjB0j6/e2LrH9xfOFtyEDqccBDaUXUQiqeC/sxzDSAIAYIQiEFikBgjBolBYpAYJAaJQRmOQYIQlDItNHXNv/3uaG7ZIHQ44SC0o+ogZCoIQBACBCEQg8QgMUgMEoPEIDFIDBKDmiEGCUJQutv3Ta77g/uHzy4YhA4nHIR2VBWETAUBCEKAICQIIQaJQWKQGCQGiUFikBgkBjVTDBKEoDwbD0yt+otHR082NAjtqCoImQoCEIQABCHEIDFIDBKDxCAxSAwSg8SgZotBghBU5o7HJ9f80bcKM4kHoR0VByFTQQCCEIAghBgkBolBYpAYJAaJQWKQGNSsMUgQgmqmhSZX3bh17PCTe29NJgjtqDgImQoCEIQABCHEIDFIDBKDxCAxSAwSg8SgZo5BghBUr/Pop1+vexDaUb6N39v6G1NBAIIQgCCEGCQGiUFikBgkBolBYpAYJAYJQlAD//knK/fVNQjtqMzY0f/xq54fAEEIQBBCDBKDxCAxSAwSg8QgMUgMEoMEIUh7ENpRuf/843/5V54fAEEIQBBCDBKDxCAxSAwSg8QgMUgMEoPOBaEpQQhSGYR2CEIAghCAIIQYhBgkBiEGiUFikBgkBglCkN0gtEMQAhCEAAQhxCDEIDEIMUgMEoPEIDFIEILsBqEdghCAIAQgCCEGIQaJQYhBYpAYJAaJQYIQZDcI7RCEAAQhAEEIMQgxSAxCDBKDxCAxSAwShCC7QWiHIAQgCAEIQohBiEFiEGKQGCQGiUFikCAE2Q1ChwQhAEEIQBBCDEIMEoMQg8QgMUgMEoMEIchuEDpUjyC0QhACEIQABCHEIDEIMUgMEoPEIDFIDBKD5gehaUEIGhWEDtUjCK0QhAAEIQBBCDFIDEIMEoPEIDFIDBKDxCBBCFIRhA7VIwitEIQABCEAQQgxSAxCDBKDxCAxSAwSg8QgQQhSEYQO1SMIrbg0CP1IEAIQhAAEIcQgMQgxSAwSg8QgMUgMEoMEIahREPrv91Ubg6oPQisEIQBBCEAQQgwSgxCDxCAxSAwSg8QgMWhh44IQJBuEDtUjCK0QhAAEIQBBCDFIDEIMEoPEIDFIDBKDxKDFY5AgBAkGoUP1CEIrBCEAQQhAEEIMEoMQg8QgMUgMEoPEIDFo6RgkCEFCQehQPYLQCkEIQBACEIQQg8QgxCAxSAwSg8QgMUgMWj4GCUKQQBA6VI8gtKKEIPQvBCEAQQhAEBKDxCAxCDFIDBKDxCAxSAwSgwQhqHsQOlSPILRCEAIQhAAEIcQgMQgxSAwSg8QgMUgMEoNKj0GCENQxCB2qRxBaIQgBCEIAghBikBiEGCQGiUFikBgkBolB5cUgQQjqFIQO1SMIrRCEAAQhAEEIMUgMQgwSg8QgMUgMEoPEoPJjkCAEdQhCh+oRhFYIQgCCEIAghBgkBiEGiUFikBgkBolBYlBlMUgQghoHoUP1CEIrKvKPB//rH3t+AAQhAEFIDEIMQgwSg8QgMUgMEoPEIEEIahmEDtUjCK0QhAAEIQBBCDFIDEIMEoPEIDFIDBKDxKDqYpAgBDUKQofqEYRWCEIAghCAIIQYJAYhBolBYpAYJAaJQWJQ9TFIEIIaBKH/WI8gtEIQAhCEAAQhxCAxCDFIDBKDxCAxSAwSg2oTgwQhSGMQWiEIAQhCAIIQYpAYhBgkBolBYpAYJAaJQbWLQYIQ1CII/Xc1DEIrBCEAQQhAEEIMEoMQg8QgMUgMEoPEIDGotjFIEII0BaEVghCAIAQgCCEGiUGIQWKQGCQGiUFikBhU+xg0PiEIQTqC0FV1CEL/lSAEIAgBCEJiEGIQYpAYJAaJQWKQGCQGCUKQjiB0lSAEIAgBCEKIQWIQYpAYJAaJQWKQGCQG1S8GCULQ6CB0lSAEIAgBCEKIQWIQYpAYJAaJQWKQGCQG1TcGCULQyCB0lSAEIAgBCEKIQWIQYpAYJAaJQWKQGCQG1T8GCULQqCB0lSAEIAgBCEKIQWIQYpAYJAaJQWKQGCQGJRODBCFoRBC6ShACEIQABCHEIDEIMUgMEoPEIDFIDBKDkotBghAkHYSuEoQABCEAQQgxSAxCDBKDxCAxSAwSg8SgZGOQIARJBqGrBCEAQQhAEEIMEoMQg8QgMUgMEoPEIDEo+RgkCEFSQegqQQhAEAIQhBCDxCDEIDFIDBKDxCAxSAxqTAwShCCJIHSVIAQgCAEIQohBYhBikBgkBolBYpAYJAY1LgYJQlDvIHSVIAQgCAEIQohBYhBikBgkBolBYpAYJAY1NgYJQlDPIHSVIAQgCAEIQohBYhBikBgkBolBYpAYJAY1PgYJQlCvIHSVIAQgCAEIQohBYhBikBgkBolBYpAYJAalIwYJQlCPIHSVIAQgCAEIQohBYhBikBgkBolBYpAYJAalJwYJQlDrIFRZDPrHg/UIQv+lIAQgCAEIQmIQYpAYJAaJQWKQGCQGiUFikCAEtQlCv7Wv2hgkCAEIQgCCkBiEGIQYJAaJQWKQGCQGiUF1i0GCENQqCFUXgwQhAEEIQBASgxCDEIPEIDFIDBKDxCAxqG4xSBCCBgahg4IQgCAEIAiJQYhBiEFikBgkBolBYpAYlEAMEoSgQUHoYAJBqEUQAhCEAAQhMQgxSAwSg8QgMUgMEoPEIDFo1qQgBEkHoYMJBKHtghCAIAQgCIlBiEFikBgkBolBYpAYJAaJQedjkCAECQehgwkEoe2CEIAgBCAIiUGIQWKQGCQGiUFikBgkBolB82JQbEIQgmSC0MEEgtB2QQhAEAIQhMQgxCAxSAwSg8QgMUgMEoPEoMtikCAECQWhgwkEoe2CEIAgBCAIiUGIQWKQGCQGiUFikBgkBolBC8QgQQgSCEIHEwhC2wUhAEEIQBASgxCDxCAxSAwSg8QgMUgMEoMWiUGCENQiCP3LfdXGoKqC0HZBCEAQAhCExCDEIDFIDBKDxCAxSAwSg8SgJWKQIAR1DEIHEwhC2wUhAEEIQBASgxCDxCAxSAwSg8QgMUgMEoOWiUGCENQpCB1MIAhtF4QABCEAQUgMQgwSg8QgMUgMEoPEIDFIDCohBglCUIcgdDCBILRdEAIQhAAEITEIMUgMEoPEIDFIDBKDxCAxqMQYJAhBjYPQwQSC0HZBCEAQAhCExCDEIDFIDBKDxCAxSAwSg8SgMmKQIAQ1DEIHEwhC2wUhAEEIQBASgxCDxCAxSAwSg8QgMUgMEoPKjEGCENQoCB1MIAhtF4QABCEAQUgMQgwSg8QgMUgMEoPEIDFIDKogBglCUIMg9OMEgtB2QQhAEAIQhMQgxCAxSAwSg8QgMUgMEoPEoApjkCAEAQSh7YIQgCAEIAiJQYhBYpAYJAaJQWKQGCQGiUFVxCBBCFIehLYLQgCCECwgPzy6BaoxMjp+aGx8KqIak6TY6HxjZM8E540sZpT6Gi9bHAHEIDFIDBKDGhmDBCFIcRDaLggBCEKwiIHBQgQAQDjizWwxSAwSg8SgRsYgQQhSGoS2V+//e+6f9Xl+AAQhBCEAAAQhMUgMEoPEoHNBaFIQglQFoe01CkIH/tmo5wdAEEIQAgBAEBKDxCAxSAwShCBtQWi7IAQgCIEgBAAgCIlBYpAYJAbVOAYJQlCLIPQvahOEtgtCAIIQCEIAAIKQGCQGiUFiUB1ikCAEKQlCLYIQgCAEghAAgCAkBolBYpAYVKcYJAhBCoJQiyAEIAiBIAQAIAiJQWKQGCQG1TEGxYrP72pramhQEGoRhAAEIajA4NDICRsrAACCkBgkBolBYpAgBAEEoRZBCEAQgiqCUP9AIQIAIAwjo+NikBgkBolBDY1BghA0KAi1CEIAghBUHYSGIwAAwpBEEBKDxCAxSAwShCBlQahFEAIQhEAQAgAQhMQgMUgMEoMSjEGx4tf61dbUkFAQahGEAAQhqIGh/OgWGysAAOEYLoyJQWKQGCQGNTQGxaynQRACQBBCEAIAoI7yw6NikBgkBolBDY1BghAkGIRaBCEAQQhqF4Q22VgBAGjuICQGiUFikBhUpoL1NCQQhFoEIQBBCGooPzy62sYKAEA4BgYLYpAYJAaJQY2MQfFjcMJ6GuochFoEIQBBCAQhAICmJwaJQWKQGNSoGHQ+CB23noY6BqEWQQhAEII6GB4eW2lTBQAgLHFMEIPEIDFIDGpgENpiPQ11CkItghCAIAR1ZFMFACAs8YawGCQGiUFikCAEIQehf76v2hgkCAEIQlC2gcFCzsYKAEA4RscmxSAxSAwSgxqm+LWw2loaahyEWtIShP4LQQhAECLjQeiEjRUAgHCMjI6LQWKQGCQGCUKQlSDUIggBCEKQkMGhkf02VgAAwpEfHhWDxCAxSAxqGOtoqGEQahGEAAQhSNBQfmRT30A+AgAgDMX3b2KQGCQGiUGNUrCOhhoFoZYUBqGnBSEAQYiMB6HR1X39+QgAgHCIQWKQGCQGNULx8TlhHQ01CEI/SmEQ2iYIAQhCZF5+ePRqmyoAAGGJY4MYJAaJQWJQA4LQfutoyGAQ2iYIAQhCNA2bKgAAYYk3jMUgMUgMEoOSVvz62GQNDRkLQtsEIQBBiKYyMDh8wsYKAEA4RkbGxSAxSAwSgxI1di4IrbaGhgwFoW2CEIAgRPMFoaHCfhsrAADhyA+PikFikBgkBiUag2LWz5ChILRNEAIQhGhKg0Mjm2ysAACEo/j+TQwSg8QgMSjRGFT83wXrZ8hIENomCAEIQjStofzIahsrAABhEYPEIDFIDEoqBsWKj9lx62fIQBDaJggBCEI0PZsqAABhiTeSxSAxSAwSg5KIQWPjs0Foi7UzBB6EtglCAIIQFPUPDJ+wsQIAEI7RsQkxSAwSg8SgRGJQrPg1s9raGQIOQtsEIQBBCM4bGCzs7+3PRwAAhGFoeFQMEoPEIDEokRgUs26GWgah/zbZILRNEAIQhGCewaGRtb19+QgAgDD0DwyLQWKQGCQGJRKDir+Ws26GQIPQNkEIQBCCywzlR662sQIAEJY4TohBYpAYJAbVMwadvz9ov3UzBBiEtglCAIIQLKKvP1/o7RuKAAAIw+jYpBgkBolBYlBdY9D5+4PWWjNDYEFomyAEIAjBEvoHhltsrAAAhGPRe4TEIDFIDBKDahSDYsXvn5XWzBBQENomCAEIQrDcPUKDhfU2VgAAwtHfPywGiUFikBhU1xjk/iAILAhtE4QABCEo+R4hGysAACG55B4hMUgMEoPEoBrGIPcHQWBBaJsgBCAIQXn3COVsrAAAhKMwOi4GiUFikBhUlxjk/iAIKAhtE4QABCEo/x6h/TZWAADCMZgfEYPEIDFIDKpLDIpZJ0MAQWibIAQgCEEl9wgNFVbbWAEACIsYJAaJQWJQPWJQ8bE5bp0MKQ9CNYpBZwUhAEGI5tTbN3TGxgoAQDjijVsxSAwSg8SgWsag2fuDpqY3WSNDioNQDWOQIAQgCNG8x8a12FgBAAjHUMnHxolBYpAYJAaVrvg9dbU1MqQ0CL18VU1j0Ky9//Q3nh8AQYgmMzA4vL6nbzACACAMff15MUgMEoPEoJrGoOK/m7M+hpQGoZdrE4TOLsDzAyAI0XT3CI2s7OkdjAAACEe8KS0GiUFikBhUixjkuDhIcRB6uTZB6KwgBCAIwZy+/vxxGysAAOHID4+KQWKQGCQG1SQGOS4O6h2E/pt91cagaoLQWUEIQBCCK46Ns7ECABCMhY+NE4PEIDFIDCqf4+IghUHo5doEoaVi0NmtghCAIIRj4wAACMLY+JQYJAaJQWJQVTFo9ri4ScfFQaqC0Mu1CULLxSBBCEAQwrFxNlcAAAIxlB8Rg8QgMUgMqioGOS4OUhaEXq5NEColBglCAIIQzX1s3FobKwAA4ejtGxKDxCAxSAyqKgY5Lg5SFIRerk0QKjUGCUIAghBNrqd38IzNFQCAcIyMjotBYpAYJAZVc1zcemthSEEQerk2QaicGCQIAQhCODZuv40VAIBwDAwWxCAxSAwSg6o5Lm6ltTA0OAi9XJsgVG4MEoQABCGa/ti4wrU2VgAAwhJvpItBYpAYJAaVPx001WIdDA0OQi/XJghVEoMEIQBBCP5Jb99QzsYKAEA48sOjYpAYJAaJQWUrfs2ttgYmQ3/B9ZrevqGtXT0Db3R29eWW1r+07oV1XTCwsJ5zui/T2/rGB/3vvBRd4VeXeWdpA2//YEH9y7j09790iXgPaFH98+Vn9ZVi4Er9A8NVGRoaOTxcGNs8Mjpxja93QBCCGir+oF3f3TMYAQAQht6+ITFIDBKDxKCyFP/cgvUvmTj6fiC/JtfVl2tt64oW1L6Y7iu0zdexnJ4L2ufLLaf3go5ydM7pW1BuIV2L6b+gczndV+pa1MBFPVfqXlYJ73t6B6P+wUKuMDK+xtc/IAhBbf5Wzcqe3sEz3SX9sAYAIA1Gx8bFIDFIDBKDyjgubnqT9S+B712synX25U4vFoJEoUxHodjgUOHk6NjkKt8PgCAE1f4Nm/78fhsrAADhGBgcFoPEIDFIDCp1OuhM8ftupbUvAZ9scl1be/fZOAbNEYWaMwoVvxbyI6MT1/m+AAQhqOpv2gxfbWMFACAs8Sa7GCQGiUFi0PLTQVMt1r1kKQaJQs0dhXr7hs6aFAIEIahS8QfqcRsrAADhGBwqiEFikBgkBi2r+L10tTUvoR4T197RM3O6tSuaJQqJQvMmhXyPAIIQVPe3blbbWAEACEscGsQgMUgMEoOWOC7uhPUuoers7n/jdGtndCEIiUKi0LwolB8ePeD7BBCEoAo9vYMnbKwAAIQjPzwqBolBYpAYtIiJ+OtptbUuQf6l1cHha87FoDmikCh0aRRydBwgCEGV+vrz622sAACEo6c3/VNCYpAYJAY1JgaZDiIb00GikCi0eBTKD49t9f0CCEJQheIP3sJCP6wBAEinNE8JiUFikBjUmBh0fjporTUuoWpt7zp7ZRAShUShS/W5SwgQhKD6KSEbKwAA4ejpHRSDxCAxSAy6JAYV//yC9S3B7ksMDF93asEYJAqJQldybBwgCEEtpoTm/9AGACDVCiPjYpAYJAaJQRengyan11vbEuz9xn2Dm+MgJAqJQqVEoeJ7oDW+bwBBCKqdErKxAgAQjHhKKC13CYlBYpAY1NgYVPz/poMI/S+pHpgLQqKQKLRcFBKEAEEIajYltNQPcwAA0mQoBXcJiUFikBjU6BhkOojsBSFRSBRaKgoJQoAgBDWZEhpab2MFACAc8WZJI6eExCAxSAxqfAwq/jdPWM+SxSAkColCi0UhQQgQhKB2b8JyNlcAAAKaEsqPiEFikBjUpDHo/HTQamtZshqERCFRaKEoJAgBghDU7i6h1TZWAABCmhLqT3xKSAwSg8SgdMQg00E0QxAShUShy6OQIAQIQlDbN2InbK4AAIRjYHBYDBKDxKAmi0Hnp4OutYYlC7qWCUKikCg0PwoJQoAgBDXUP5C/2sYKAEBY4o1oMUgMEoOaKQZNtVi/0kxBSBQSheaikCAECEJQYz29g/sX+oEOAEA69fXnxSAxSAxqkhhU/LUzxe/LldauNFsQEoVEoZggBAhCUOu7hAbyK4s/pM/YXAEACMfI2LgYJAaJQZmPQbPTQVusW2nWICQKiUKFgiAECEJQc719Q5s6S/mBDwBAKsSbJHHEEIPEIDEouzGo+OsF61WyGYRykSgkCpUShQQhQBCCer0p6+7PdRZ/+AMAEIah/IgYJAaJQZmNQfF00PRqa1Wyt/cwF4REIVFo+Sg0LAgBghDUbUroWhsrAABhiTeNxSAxSAzKYgyaarFOJatB6P3Tc0FIFBKFlo5CghAgCEEdFX/Y7rexAgAQjr7+ITFIDBKDMhaDir/nTPH7c6U1KlkOQqKQKFRKFBKEAEEI6qivP7+y+MO5YHMFACAc+eFRMUgMEoMyE4Nmj4pbb31KMwQhUUgUWi4KCUKAIAT1PzputY0VAIBwdHX3zW72i0FikBgUfgwqfhwnrEtppiAkColCS0UhQQgQhMDRcQAAVHF0nBgkBolB6YxB8VFxxe+zq61JabYgJAqJQotFIUEIEIQgoaPjOrv6CrnF3iAAAJA6+eERMUgMEoOCjUHxUXFTm6xHyX4Q6l8wCIlCotBCUWi4MCYIAYIQJHN03OBqGysAAOGIj46LN5XFIDFIDAovBhUfp+PWoTR7EBKFRKHLo5AgBAhCkPDRcTZXAADC0dM7IAaJQWJQYDFo9qi46ZmV1qAIQqKQKHRpFBKEAEEIEtbZ1ZfLFd80AAAQhsH8iBgkBolBwcSg+Ki46bXWnjTNHkMJQUgUEoXmopAgBAhCkLCe3sFriz/sz9hcAQAIx+jYhBgkBolBAcSg4uO+37oTQUgUEoUWjkKCECAIQUOi0MB6GysAAOHo7O6b3eAXg8Qg21uQYgAAIABJREFUMSi9Maj4MeSsNxGERCFRaPEoJAgBghA07pzfFpsrAADh6OkbFIPEIDEorTEovjdoauZqa00EIVFIFFo8CglCgCAEDdLbN7TSfUIAAIHdJzRUEIPEIDEodTHIvUEIQqKQKFRKFBKEAEEIGn2fUGfvmYtvGgAASLvC6JgYJAaJQSmKQe4NoqmDUFdlQUgUas4oJAgBghA0WHfvwFobKwAA4ejs6o1GxyfEIDFIDEpDDJqYPGFdSbMHofdOdUSikChUShQShABBCNJxn9CWjnLfYAAA0DDdPf2zEUAMEoPEoMbFoOK/Uyh+/620pkQQ6ohEIVGolCgkCAGCEKQmCvW1dBTfbAAAEIbevkExSAwSgxoXg84Un7trrSWpah3eM3Bdrqtvc3uu50Bre/cbp9o6c7HTbV0VaZ2vvXRtC+peWMeliv/dmbkgJAqJQstFod6+oXxffz63oIEr9Q8MV2+wMGugHEMjs4byo2/kh8cOFArjm0dHJ67zugWCEGRGb9/gylxnb87mCgBAOPoH8mKQGCQGJR6DJuLnbq11JJWIA9Dptq6T777XfvZX77ZFV3jvnHeW1b6gd+d7v3TvLWRe6CmHKCQKlXqn0DkDF/VcqXtZg8vrPadnUUNX6ruo97y+/vzZOBIVRsbXeT0DQQgyEYWKbxjO2FwBAAhHfnhUDBKDxKBkY9B660fKuru3Z2BVPAX0znttZ3/1bmt0UVskColColBYUWhO/8DwTGFkfLPXOBCEIPQ3qtd25HpEIQCAgBRGxsQgMUgMSiAGFR//FutGytGe690ah6BfXhKCRCFRSBTKQhS6GIYmTAyBIATBRyGbKwAAgch19kajYxNikBgkBolBpOd+oGveO9WRj0PQfKKQKCQKZS8KxQbzIyfHxqdWef0DQQjCfPPa3b/e5goAQEhRqCeoKCQGiUEhxaDix5KbnJ5Zaa1ISfcEdfatm5sKWogoJAqJQtmMQv0DhZnRscnrvA6CIATBRqHl34QAAJAWcRSKN/vFIDFIDBKDaIyOzt7Nv3ynNbpAFBKFRKGmikJ9A8NnRSEQhCDkKLTJ5goAQDi6uvtSHYXEIDFIDCKzMSgXx6DT0TmikCgkColCXhdBEIIAdXb1tdhcAQAQhcQgMaipYtD45BkxiDLWzWsuxiBRSBQShUSh2Sh0jddHEIQg3ChUfIMCAEAY0haFxCAxKLQYVHz+rrUWpMSTNa751butZ68MQqKQKCQKNXMUGhgs5L1GgiAE4V6MKQoBAIhCYpAYJAbBJd4/ncstHINEIVFIFGr2KJQfHjvsdRIEIQg3CnX2ikIAAKKQGCQGiUEwe29Qz+alY5AoJAqJQs0ehdwnBIIQiEIAAGQ+ColBYpAYRNa9+377TGlBSBQShUShZo1Cg0MjOa+XIAhB4MfH9e63uQIAEI7OhKOQGCQGBRWDJiZzk9MzK631KEd7rmfzyV+VGoNEIVFIFGrmKDQyOrHG6yYIQhC0zq6+9cu/eQEAIC1ynb3R6NiEGCQGiUFiEDXwznvtM3EQEoVEIVFIFFouCg3lR9/wugmCEIhCAAAkqiPXXdcoJAaJQWIQzXFqRv91czFIFBKFRCFRqJQoVPxZtcrrJwhCkIUotLa9o/tM2+VvaAAASKU4ChVGxsQgMaipY1Dx8W+xnqNSp9u6Dl8ehEKKQn//D7+IXv3RG9G+/S/Muv/BLZf6drW+n6hv1Mt3amlrzXwzCQ/V0raKPPz9PdFTz/1d9OLLR6PX3/xpdLo1F3QUKoyMb/b6CYIQZEJXd9+1ohAAQFiGhkfEIDFIDIIKvPt+e/7kr05FoUShv/+HE9HTL7RE3350Z7Ru433Rreu/CkHa+LUHom2790cHj/34fCAKJwo5Ng4EIchWFOrpv7q9ozvX1t4VAQAQhr7+ITFIDGqqGFR87tZbv1GtczFoTjqj0GwEev7l6J7NDwkJZNbXvvFwdPDoj2aP/Et7FBoYLOS9foIgBJlS/EG6siPXc9zmCgBAOOJNijgsiEFiULZj0OSZ4nO31rqNqu8P6uxbc2kQSlcUOvbD12cngcQCmk08ORR/76U5CnkNBUEIMqmjs2e/zRUAgHB0dvXObtyLQWJQJmPQxGSu+Nxda61GTda7ud51VwahxkehYz98Ldr84BZhgKb3rYe2Ra+9+dNURqHR0YnrvI6CIATZ/FtTXb3r29q7zrS2d0UAAKRfe647KoyMiUFiUKZiUPFjOjE5PbPSGo1aKb5eHlg4CDUmCv3k9f9XCILFJobeOZ2qKDQyOrHG6ygIQpBZnV1917a1dxdssAAAhGNwqCAGiUGZiEHF522LdRnJBqHkotDPT7wT7dj7VHTLuq8Ai1i/cVP09HN/l5ooJAiBIASZ19Xdv7I913Pc5goAQDi6e/oXvFdIDBKDwohB8X1B0+4LokFBqP5R6OgPX4vuuuebNvyhRF+7/+FLpoUaFYUEIRCEoIku3uzd1NrWFQEAEIaOXE+8cSEGiUFhxaCJydzk1MzV1mDUMwj94pfLBaH6RaHH9j9vgx8qnBY6ePRHDY1CIyOCEAhC0HRHyHUVbLAAAIQjPkJODBKDQohBxcd9v3UXSQWhpKPQz068E337kZ029qFKe598vmFRSBACQQia9Qi5lta2zggAgDB0dvVFYxNTYpAYlNIYNHtE3GrrLZIOQklFoZ+9/U50933fsZkPNfLd7++NThff3yQdhQqCEAhC0MRHyK1tbes6Y4MFACAM7R1dUb4wKgaJQamKQcXH6fjk9MxKaywaFYTqHYV+fPzvozvv/oZNfKixe+//buJRSBACQQhMC3V0n7DBAgAQju6e/sWnhcQgMSixGDQ7FbTWuoo0BKF6RaE4Bt2x4Ws27yEjUUgQAkEIKOro7Fnf2tZpWggAIBBtC00LiUFiUEIxyFQQaQxCtY5CP3v7V46Jg4SiUFJ3ChVGxgUhEISAWGd3XzwtdDz+mxkAAIQhnhYaHZ8Qg8SghGKQqSDSHYRqFYXEIEjW1l1PJhKFBCEQhIArp4XWtrZ1FmywAACEoa29KxoYHBaDxKC6xqDi87R/ylQQAQShWkShR7bujW5Z92UgQU89+1Ldo5AgBIIQsNC0UNfstNCW062dEQAAYejo7ImGC2NikBhU0xhU/O/nil8jq62TSIvTbcsHoWqi0P5nXoq+cMeXgQZ47c2f1jUKCUIgCAFLh6Gr29q7TpxuzUUAAIQh3iQZHZsQg8SgKmPQ7PFw662LSGcQej+qRxT60U/+3qY8NNC6u74+O/1crygkCIEgBJRyjFyuZ/XsMXI2WAAAgtDW3hn19Q9FY+NTYpAYVHYMcjwcYQSh2keh+N4gm/LQWN/dsudCEKp1FBKEQBACygtD60+3dp6xyQIAEEgY6uiOhvIFMUgMKikGFZ+blsmpmautfQgnCNUuCu154jmb8ZASP/zxG3WJQoIQCEJA5fcLCUMAAMGGITFIDLrknqAT7gki3CBUfRR6/a2f2YSHFNlw9zcvOTquVlFIEAJBCBCGAACaRq6zLxoujIhBYpAQRMaCUHVR6IGHt9uEh5R56tmXLglCtYhCghAIQkANwlDbbBjKnTnVmosAAEi/XGdPNDhUEIOaNAYJQYQehE4sGIQqi0JHX/2JzXdIoTvu/NoVU0LVRiFBCAQhQBgCAGhabe1diYQhMSgdMWg2BE0JQWQjCNUqCn3ru6aDILVTQs9cOSVUTRQShEAQAmos19UbHyW3/nRrrnDqdC4CACD94jDU2zc0Gw7EoOzFoOLz0DI5PXO19QpZC0LVRqFzdwdtBFIqnhLq6h6oWRQShEAQAuqovaN7bWtb5wmbLAAAYWhty0VdPf3R6Ni4GBR4DCr+2WeKz8EWIYisB6FqotDD399j0x1SruXIf6hZFBKEQBACkpga6uy9urW9q+VUfJycjRYAgCBUe8+QGNSYGFT8nOP7gdZbh9BMQajSKPSlO++NPv+ljUCK3bP5oXNBqAZRSBACQQhINgzNHSeXO3W6IwIAIP3iqaGe3sGypobEoGRj0PlpoP1TpoFo4iBUbhR69m8P2WyHQMTfs7WIQoIQCEJAg3Scmxraf6o1V3j/dEcEAED6tXd0R/0D+SXvGhKDkotBxc/z+OTU9FrrCwSh8qPQtx7aZqMdAvH8S4cvBqEqopAgBIIQkI67hq5tbetsOXW644yNFgCAMHR29UWDQ8OXxCExqP4xKI5A8ZFwU9MzK60laMog1Nq5ZBAqNQrZZIdw3H3fd6Ku7v6qo5AgBIIQkL44tLq1rXP/qdMdJocAAAKKQ30DQ9HI2LgYVIcYVHyMjk9MiUBwIQidXDoILReFDh/7jzbZITCnWnNVR6FCQRACQQhIrbZzk0Nbij/0czZaAADC0NbRFXX3DkT5wogYVGEMKv7+wsTkVEt8HJwIBIsEoSqi0O59z9hgh8C8+h9eOx+EKo9CghAIQkAwdw71rGzr6F57/mi5wvunOiIAANIt/tu8ua7e2emh4ZExMWiJGDQxOXsf0Kaia73/hxKDUIVR6OvfeMQGOwRm9+PPzAtClUWhYUEIBCEg0ECU67m6rb1r/fnj5XLvn2qPAABIt1OtHbOBqLdvMMoPjzRtDCr+8zNxACraMjk1vdr7e6giCFUQhT7/xY1AYO5/cMtlQaj8KCQIgSAEZOuIufj+oS2nW3PHz00R2XQBAEi71vauqKu7L+rrH5qNRKNjk5mKQXH8GZ+cOjExObV/8tw9QFd77w41DkJlRKHX3vypzXUI0Jf+5t4FglB5UUgQAkEIyHokau9afX6SKA5FJ0wTAQAEEInaOqOOXPfs5s1cKBoujKU9BsVTP3H4aZmb/BF/oPZOLRaESoxCh4/9OPrLL94FBGjhIFR6FBKEQBACmvvIuYuxqK1zfxyMYu+bLgIASO+xc6c7ZmNRrKdvYNZcNJozOjZR8+BzPvacmDvqbS76OPINkg9Cby8WhEqIQk88/bc21iFQP3n9P1UVhQQhEIQASp0yWsza0+eCElSlu3fgpz19g7+si97lDABp03NOd0X6ocb6Uq2rAkPDo387OTW9aS7oLMR0D6Q7CFUahXbue8bGOgQchDoXDULLRyFBCAQhAAAAAAIMQpVEIUEIwvXy4R/OBqFKo9BwYUwQAkEIAAAAgHCC0HtRpVFoy47HbaxDoJ448OKFIFRJFBKEQBACAAAAILggVFkUuvf+79pYh4wEoXKjkCAEghAAAAAAQQah8qOQIAQBB6GnrwxC5UQhQQgEIQAAAACCDULlRSFBCAIPQl39FUchQQgEIQAAAACCDkKlR6HZIHT7BiBAF4JQhVFIEAJBCAAAAICQgtAvFgpCpUWhOAjdfPsGIECXBKEKopAgBIIQAAAAAKEFoQqjkCAEGQpCZUYhQQgEIQAAAACCCUK5i0GogigkCEHGglAZUUgQAkEIAAAAgFCDUJlRSBCCDAahEqOQIASCEAAAAAAhB6EyopAgBOF6fKkgVEIUEoRAEAIAAAAgEO8vFoRKjEKCEAQchJ5aJggtE4UEIRCEAAAAAMhCECohCt0jCEHQQSi3XBBaIgoJQiAIAQAAABBKEDq9TBBaJgoJQhB+EKo0CglCIAgBAAAAkKUgtEQUumfzQ9HNt98JBOjxp164EIQqiUL5YUEIBCEAAAAAshWEFolCs0HotjuBAJ0LQn0VRyFBCAQhAAAAALIYhH6xcBC66bY7gQBdDEKVRaH88KggBIIQAAAAAKEEoZ//4t2o0igkCEFWglD5UUgQAkEIAAAAgMCCUKVRSBCCLAWh8qKQIASCEAAAAAABBqFKopAgBFkLQqVHIUEIBCEAAAAAQgpCJy4GoXKjkCAEWQxCpUUhQQgEIQAAAABCC0IVRiFBCMK1Lw5CnX0VRyFBCAQhAAAAAEIMQhVEIUEIMhCEKoxCghAIQgAAAACEGoTKjEKCEGQkCFUQhQQhEIQAAAAACDkIlRGF7r7voeimW+8EArRv/2VBqMwoJAiBIAQAAABA6EGoxCh0933fiT53698AAXpsoSBURhQShEAQAgAAACALQaiEKCQIQdhBqGOhIFRiFBKEQBACAAAAIJQgdGqZILRMFBKEIPwgVGkUGsoLQiAIAQAAAJCdILREFBKEIOQg9PyFIFRJFBKEQBACAAAAIGtBaJEoJAhBdoJQuVFIEAJBCAAAAIBAvHeqo/QgtEAUEoQgW0GonCgkCIEgBAAAAEBAQehnJ96JKo1CX90kCEHWglCpUUgQAkEIAAAAgMCCUKVRSBCC0INQb8VRSBACQQgAAACAAINQJVFIEIKAg9CTc0GosigkCIEgBAAAAECgQajcKPTVTd+O/v0tfw0EaG8chHK9FUchQQgEIQAAAAACDkLlRCFBCDIQhCqMQoIQCEIAAAAAhBSE3r4yCJUahQQhyEgQqiAKCUIgCAEAAAAQWhCqMAoJQpChIFRmFBKEQBACAAAAIMQgVEEUEoQg4CD0xAJBqIwoNJQfEYRAEAIAAAAgyCBUZhQShCCDQajEKCQIgSAEAAAAQMhBqIwoJAhBRoNQCVFIEAJBCAAAAIDQg1CJUUgQgpCD0HNLB6FlopAgBIIQAAAAAFkIQiVEoa/MBqG/AgJUUhBaIgoJQiAIAQAAABCId5cLQstEIUEImiAILRKFBCEQhAAAAAAIKAj9dLkgtEQU+srXH4w++4W/AgJUVhBaIAoJQiAIAQAAABBYEKo0CglCEHYQai8nCF0WhQQhEIQAAAAACCYItV8IQpVEoa98/QEb6xCoPeeDUKVRSBACQQgAAACAoILQr6JKo5AgBCEHoWcvBKFKotCgIASCEAAAAAChBaHKopAgBKEHoZ6Ko5AgBIIQAAAAAEEGofKjkCAEAQehx+eCUGVRaHBIEAJBCAAAAIBAg1B5UUgQgqwEofKjkCAEghAAAAAAQQeh0qPQV772QPTZz68HAnRlECovCglCIAgBAAAAEHwQKi0KCUKQtSBUehQShEAQAgAAACATQWj5KCQIQRaDUGlRSBACQQgAAACAUILQ+8sFoaWj0Je/9kC09vPrgQDtefyZJYLQ8lFIEAJBCAAAAICQgtDPlwtCi0ehL98rCEF2g9DSUUgQAkEIAAAAgNCCUIVRSBCCwINQR0/FUUgQAkEIAAAAgBCDUAVR6Mv3fsvGOoQehCqMQoIQCEIAAAAAhBqEyoxCghCEa/f8IFRBFBKEQBACAAAAIOQgVEYU2igIQbB2Pf5M1DY/CJUZhQQhEIQAAAAACD0IlRiFBCEIPwhVGoUEIRCEAAAAAMhCECohCs0Gob9cDwRo176LQaiSKCQIgSAEAAAAQFaC0M9LCULrgACdC0LdFUchQQgEIQAAAACyFISWiEJ33fut6Ma/XAcE6GIQqiwKDQ4VBCEQhAAAAAAIJwj9Mqo0Ct11jyAE2QhC5UchQQgEIQAAAACCC0KVRSFBCLIUhMqLQoIQCEIAAAAABBSE/uFCECo/CglCkLUgVHoUEoRAEAIAAAAgsCBUaRS6655v2liHYIPQgUWCUGlRSBACQQgAAACAAINQJVFIEIKsBqHlo5AgBIIQAAAAAIEGoXKjkCAEAQehx5YLQktHoQFBCAQhAAAAAMINQuVEIUEIAg9C7d0VRyFBCAQhAAAAAALxznttCwahUqPQbBC6+Q4gQDvnglCFUWhgUBACQQgAAACAcILQzxYOQqVEoTgI3XDzHUCALglCFUQhQQgEIQAAAABCC0IVRiFBCMIOQq3zg1CZUUgQAkEIAAAAgBCDUAVRaIMgBMEHoUqjkCAEghAAAAAAoQahMqPQhrsFIQg2CO29GIQqiUKCEAhCAAAAAIQchMqIQoIQZCcIlRuFBCEQhAAAAAAIPQiVGIU23P0NG+sQbBB6+oogVE4UEoRAEAIAAAAgC0GohCgkCEHoQair4igkCIEgBAAAAEBWgtAyUUgQgiwEocqikCAEghAAAAAAAQWh/7RcEFoiCs0GoZu+BARo596n5gWh8qOQIASCEAAAAACBBaFKo5AgBFkKQuVFIUEIBCEAAAAAAgxClUShOAituelLQIAWDkKlRyFBCAQhKvdbRf9/e/cdJnddJ3D8OQvFioi9FwQbqNe9ljvvvH6nIhpRQRAU5Q7QQxA90FNBRDlUyvGgQhJI7z2bbC/JbuomW7LZlkZP3d6SzGVmdjZtZqdukt/kled5PU+e5I95dvY339/n+30/MzMuaA4d79DxDgXewXgOpuPgKXFgNAdy4UBWhlIxNJaG4hpMx+DYGxgcTN3A2OlPaiC+/uz1ZauvPyu9udAbT9+oenKpJ1W947pzqTs1XSfoyU5XYp1p605d5xEdOdWVWEfXuP1jrjNqf+e4fSdJ+LFGHneMfq6OoyV8jrP73XXGk/I1lfp1mvCaz/h1dOLrMulrOQdrRs+IJGtVlmti4rU3zlqd4bqf0T0nzftbVvfXY+7Xo9/js5ohks4vQxE5mZuSzG3xZ78M58hR5tfUZuE0Zu44s3z2e4UE+5aj9jtjt78a3icO7x/T3H86NzhJQSjdKCQIQT4GodSikCAEghCZCw+4gftz6HiHjnco8A7GczAdB0+JA6M5kAsHsjKUiqGxNBTXYDoGx97A4GDqBsZOf1ID8fVnry9bff1Z6c2F3nj6RtWTSz2p6g1151J3arpO0JOdrsQ609adus4jOnKqK7GOrtD+MdcZtb8ztO8kCT/WyOOO0c/VcbSEz3F2v7vOeFK+plK/ThNe8xm/jk58XSZ9LedgzegZkWStynJNTLz2xlmrM1z3M7rnpHl/y+r+esz9evR7fFYzRNL5ZSgiJ3NTkrkt/uyX4Rw5yvya2iycxswdZ5bPfq+QYN9y1H5n7PZXw/vE4f1jmn+cG5zEIJROFBKEILh+HQ5CDc0ZRyFBCAQhBCFBSBAShAQhQUgQEoQEIUFIEBKEBCFBSBAShAJiXW193CCUahS6WRCC4AehDKPQtu1PCUIgCCEICUKCkCAkCAlCgpAgJAgJQoKQICQICUKCkCAUmCBUtSaUaRQShCBPglAGUUgQAkEIQUgQEoQEIUFIEBKEBCFBSBAShAQhQUgQEoQEoaAFoQyj0M23CkIQ2CD08HFBKM0oJAiBIIQgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgJQoJQEINQBlFIEII8C0JpRKGtghAIQghCgpAgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgFNAilGYUEIcjDIJRiFBKEQBBCEBKEBCFBSBAShAQhQUgQEoQEIUFIEBKEBCFBKChBaEOcIJRGFLr51h+Exl95PRBAowahFKLQ1m2CEAhCCEKCkCAkCAlCgpAgJAgJQoKQICQICUKCkCAkCAUmCJXHC0IpRqFwEPr8ldcDAfSrZEEoSRQShEAQQhAShAQhQUgQEoQEIUFIEBKEBCFBSBAShAQhQShgQSjTKCQIQbCDUF2yIDRKFBKEQBBCEBKEBCFBSBAShAQhQUgQEoQEIUFIEBKEBCFBKIBBKJModJMgBAEOQr+LBKFMo5AgBIIQgpAgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgJQgENQulGIUEI8iMIZRKFBCEQhBCEBCFBSBAShAQhQUgQEoQEIUFIEBKEBCFBSBAKcBBKJwrd9B1BCPIlCKUbhQQhEIQQhAQhQUgQEoQEIUFIEBKEBCFBSBAShAQhQUgQCngQSjUKCUIQ4CD00IlBKJ0oJAiBIIQgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgJQoJQHgShVKLQTd+508E6BNQvw0GovjnjKCQIgSCEICQICUKCkCAkCAlCgpAgJAgJQoKQICQICUKCUJ4EoWRRSBCCPAhCGUYhQQgEIQQhQUgQEoQEIUFIEBKEBCFBSBAShAQhQUgQEoTyKAiNFoWiQejrQAAdE4QyiEKCEAhCCEKCkCAkCAlCgpAgJAgJQoKQICQICUKCkCAkCOVZEEoUhcJB6HNf/joQQNEgtCXjKCQIgSCEICQICUKCkCAkCAlCgpAgJAgJQoKQICQICUKCUB4GoXJBCPIrCD0YC0KZRaH2bTsFIRCEEIQEIUFIEBKEBCFBSBAShAQhQUgQEoQEIUFIEApOEFodyjQKCUKQL0Eo/SgkCIEghCAkCAlCgpAgJAgJQoKQICQICUKCkCAkCAlCglDgglBmUUgQgnwKQulFIUEIBCEEIUFIEBKEBCFBSBAShAQhQUgQEoQEIUFIEBKEAmLtMUEo/Sh0oyAEeRaEUo9CghAIQghCgpAgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgFKAiVHROE0otCN94iCEH+BaHUopAgBIIQgpAgJAgJQoKQICQICUKCkCAkCAlCgpAgJAgJQgELQplGIUEIgh2ENiUMQsmjkCAEghCCkCAkCAlCgpAgJAgJQoKQICQICUKCkCAkCAlCQQlC648EoUyiUDQIfQ0IoF8++NtIEMo0CrVvFYRAECJT5w1HoUA5dLxDxzsUeAfjOZiOg6fEgdEcyIUDWRlKxdBYGoprMB2DY29gcDB1A2OnP6mB+Pqz15etvv6s9OZCbzx9o+rJpZ5U9Y7rzqXu1HSdoCc7XYl1pq07dZ1HdORUV2IdXeP2j7nOqP2d4/adJOHHGnncMfq5Oo6W8DnO7nfXGU/K11Tq12nCaz7j19GJr8ukr+UcrBk9I5KsVVmuiYnX3jhrdYbrfkb3nDTvb1ndX4+5X49+j89qhkg6vwxF5GRuSjK3xZ/9MpwjR5lfU5uF05i548zy2e8VEuxbjtrvjN3+anifOLx/THP/6dxgLINQ5ZEglG4UEoQguO4/KghlEoUEIRCEAAAAAAhMEKqLBqEMo5AgBPkThNKNQoIQCEIAAAAABDEIZRCFbrzljtDlX/oaEEDxglA6UUgQAkEIAAAAgKAGoTSjkCAE+ReEUo1CghDKlALPAAASXUlEQVQIQgAAAAAEOQilEYXuue9hB+uQh0EolSgkCIEgBAAAAEDQg1CKUUgQguCaOnPBqEEoWRQShEAQAgAAACAfglAKUeie+x5ysA4BNXdhQdIgNFoUEoRAEAIAAAAgX4JQkij00KOTHKxDngehTYIQCEIAAAAAnAFBaJQo9OS0uQ7WIaA21TelHIQ2CUIgCAEAAABwBgShBFFoeVFF6PIvXgcEzDXXf3s4CGUehQQhEIQAAAAACIg16QShBFHoiqtvcMAOAXPzrT8MbaxryioKCUIgCAEAAAAQqCBUE8omCt1y+48csEPA/O8Dv4kEoWyikCAEghAAAAAAgQtCmUehn973YOizX7wOCJA5CwpGglCmUUgQAkEIAAAAgCAFoYpYEMosCs2Ys9gBOwTM0TEo0yjUJgiBIAQAAABAwIJQllEo/D1CDtkhGG674+64QSjdKCQIgSAEAAAAQGCC0KYjQSiLKHT7D+9x0A4B8dCjkxIGoXSiUNvWHYIQCEIAAAAABDIIZRiFfjNhmoN2CIjqNbWjBqFUo5AgBIIQAAAAAEEOQhlGoau+drPDdjjN3XrHXUljUKpRSBACQQgAAACAoAShdQmCUAZR6O6fP+jAHU5zk2fMTzkIJYtCghAIQgAAAAAEKAiVJgpCaUahgqKK0GevuBY4TV399W+lFYOSRSFBCAQhAAAAAAIWhHIVhW6/8x4H73Ca+t3E6RkFoURRSBACQQgAAACAAAahXEShBYsLQ5ddcS1wmgm/O6h20+aIXEUhQQgEIQAAAAACGoRyEYV+cNd9DuDhNPO7idNGglCuopAgBIIQAAAAAAEOQtlGofB3CX3hK990CA+niRu/c+cxMShXUUgQAkEIAAAAgEAFoepQrqPQg49MdBAPp4klBSVxg1C2UUgQAkEIAAAAgMAFodxHoRu+9X2H8XCK3ferRxPGoGyjkCAEghAAAAAAgQxCuY1CCxYXhsZf9Q2H8nCKXH/jbUljUDZRqK1dEAJBCAAAAIDgBKHyo4NQbqPQoxOmOpiHUyD8PV6LR/mouFxEIUEIBCEAAAAAghaExjAK3XXvA6HLrvgqcBL9duK0tGJQJlFIEAJBCAAAAIAgBqExjELfveOnocu+8FXgJPjFrx4J1W5szCgIpROFBCEQhAAAAAAIahAaoyhUUFQRuu6GW0Kf+cJXgTH03z+6NxqDYsYwCglCIAgBAABAWg4dOvR7MQcPHnrRwYMHRxw4cODFMUNDQy+JGRwceung4OBLBwYGz4oaOKu/f+DsqP6z+/r7z4no6zunt6/v3N7e3oie3t6X9fT0RHT39Ly8u7vn5V3d3a+I6Op+RWdX1ysjOrte2dHZ+aqIjs5X7+/oePX+/R3nhe3bt/+8vfv2vyZi777X7Nm77/yIPXvP371n72t3794TsWv3ngt27dod8cKu3a974YVdr39+2HPPv/CGmGefe/6NMc88+9ybwp5+5tk3Rzz9zFueGrbzqaffGrNj51NvC9u+Y+fbh71j2/YdEVu373jn1m3b39m+dfu7ora9q61927ujtr6ntS2qpa39vS2t7e9tbm27MKKl9cItza3vi2q5qGlLy0WbtzRfHNHUfHFj05b3R2ze8oGGxqaYD9Y3bP5gXcPmD0XUN354U31DVF3DJRvr6iNqN9VfWrux7tING+s+ElG76aPrh63bsPFjYWvX1/5+xLoNf7AmZu36P1w9rGbNuj867I+rV6+Nqln7J6tq1kSsrF79p4d9PKxqVc3Hq1bW/FnlyuqIiqrqP6+oWvUXYeWVYSv/sqyiKqK0vOqvSssrx4WVlFWOKy6r+OuI0oq/KSopP6zsE2GFxWWfWFFc+rcRRaV/t7ywJOaTBSuKP7lsRfHfRywv+oelywujCgr/ccmyFf+0OGbp8n9eNGzhkoJ/Wbh42b+GLQhbtPTf5g+bt3DJv89bsORTYXMXLP7U3PmLPh02Z/6iz8yet/Azs+cuvCxs1twFl82cM/+zwy6fMXve5TNmzftc2PRZcz8/bWbMnPFTZ8yOmDJ99hemTJ91xeRpMTO/WFq+qvyEICQKQX7EoDGOQoIQCEIAAAAgCAlCglDQg9AYRqFrRSHIfQz6n3tDGzY2RpysKCQIgSAEAAAAgpAgJAgFKAiVJApCYxiFvnvH3Q7xIUd+/stHRmLQyYxCghAIQgAAACAICUKCUMCC0MmOQmF33fuAw3zIwvirvhH6zeNTT4hBJysKCUIgCAEAAIAgJAgJQgEMQqciCj36+NTQ56+83uE+pOmq624OLVpanDAGnYwo1CoIgSAEAAAAgpAgJAgFMwidiii0YHFh6Js3f88hP6ToJ/f8KrSyZn3SGDTWUUgQAkEIAAAABCFBSBAKcBA6FVEo7IFHJkTfLTT+GiCOq667KTRrzpLQhtrGqI2NpzQKCUIgCAEAAIAgJAgJQgEPQqcqChUUVYTu/PEvHP7DUcLfFfTz+x8Jra9tjNhwtFMYhQQhEIQAAABAEBKEBKGABKGCwtIHEwWhUxWFwuYvLgzd9t93hz49/ho4Y4VD0L33PxKqrF4/EoNOpyjUvnXnJeYYEIQAAABAEBKEBKEgBKEVowehUxmFYmHoJ/f+OvTla/9TIOCMcdV1N4YefXxqqLJ6XWh9bcMJMeh0iUJmGBCEAAAAQBAShAShgAShJ6fO/FJJ2ehB6FRHoZhHH58Suu2OuyPfMyQakI8R6Ef3/DK0cEnRcAQ63ukVheobW3aaYUAQAgAAAEFIEBKEAhSEyipqnglKFCqripo+Z1Hornt/Hfrmzd8TiAhsAPqv238U+vXDj0ci0Lq4Eej0jUJNze1zzTAgCAEAAIAgJAgJQoF6h9DKZZEgFLAoFFY+bHlRRWjS1DmhBx6ZELrr3gci7vzxLyLBKN/ckMy3iPh2Mt8/KX52/8MjJk2eHZoxe3GoctW60LoNDceqbQhUFGpp236DGQYEIQAAABCEBCFBKEBBaMHigttHglCAo1DUmpRVxLNybVyVyayKr2rEuuSqk1k/YmUyNSdaVbMhdauPqF5dm7o18WwcUZPI2tGtjmtTUmvWJVN3grXr01F/xIb41sXVEF9AotDGuqY+8wsIQgAAACAICUKCUMCCUFhp7GPjRCFRSBQShZJEIR8XB4IQAAAACEKCkCAU0CBUVFo165ggJAqJQqKQKJQgCrVt3XGJ+QUEIQAAABCEBCFBKIBB6IkpM75UWlG9RxQShUQhUWi0KLS5qa3Y7AKCEAAAAAhCgpAgFOAgVLCi5KETgpAoJAqJQqLQcBQKf3eQdweBIAQAAACCkCAkCAU8CD0xZfqXS8ur14pCopAoJArFi0LNLVvvN7eAIAQAAACCkCAkCOVBEJo1Z8F/xP3oOFFIFBKFzugo1Li5dY2ZBQQhAAAAEIQEIUEoT4JQ2KJlhfeUVNQMikKikCgkCoVjUH1D8862rTvfYGYBQQgAAAAEIUFIEMqjIDRp8vQrFy1bIQqJQqKQKBSqE4NAEAIAAABBSBAShPI3CE2cPO3KRUtX/EwUEoVEoTM3ColBIAgBAACAICQICUJnQBCa+OS0q8JRqLSiZq8oJAqJQmdWFKpvbG5qa98hBoEgBAAAAIKQICQInQlBKGz6rHk3FpetXCcKiUKi0JkRhZq2tE8wn4AgBAAAAIKQICQInWFBaMITUw+b8pWly4v+ryzeu4VEIVFIFMqLKBR+V1Br+/ZLzCYgCAEAAIAgJAgJQmdwEAp7fNKUq1cUlc8tLa9+VhQShUSh/IhCDY0ta1pat403k4AgBAAAAIKQICQICUIjQeixSZOvfmzi5Gtmz1v0g8LiihUlsTgkColColBgolB9Y8uapub2+1vbvCMIBCEAAAA4NUHosIMjDhw48KKYoaGhEYODQy8eHBx88cBAzMCL+/sHXhLV/5K+mL6+l/T29b20t7c3oiespyeiu6fnrO7unrO6urujurrP6uzqOjuis+vsjs7OqI7Oc/Z3dJyzf3/Uvn37z9m7b/+5EXv3nbsnZs/ec3fv2fuy3bv3ROwK27U74oVdu1/+wgu7Xv78sOeef+EVMc8+9/yIZ5597pVhTz/zbNTTz7zqqWE7n3p6xI6dT706bPuOnTHnbdu+I2Jr2Lbt57Vv3f6aqG2vaWuP2Xp+a1tUS1v7+S2t7ec3t7a9NqKl9bVbmmNaLmja0nLB5i3NUU3NFzQ2bXldxOYtr2tobIp5fX3D5tfXxdQ3vmFTfUNUXcMbNtbVR9Ruqn9j7ca6N26Iqd30pvXD1m3YGLF2fe2bI9ZtePOamLXr37J6WM2adWFvrV69Nqpm7VtX1ayJWFm9+m0xVatq3la1subtlSurIyqqwla9I6y8MmzlO8oqqiJKy6veWVpeGVFSVvnO4rKKd0WUVryrqKT8sLJ3hxUWl717RXFpVFHpe5YXlowoWFH8nmUrit8bsbzovUuXF0YVFF64ZNmKCxfHLF3+vkXDFi4peN/CxcsuClsQtmjpRfOHzVu45OJ5C6LmLlh88dz5i94fNuew2fMWvn/23IUfCJs1d8EHZs6ZH/PBGbPnfXDGrKjps+Z+aNrMmDkfmjpjdsSU6bM/PGX6rA9PnhYz85Inp0Y9MWXGYdMvDZs0efqlEydPu3Tik9M+EjbhiamHTYl4fNKUjz42afJHH5sY9bsJT37st8OKy6q+W1qx6p7ylWsWhlUcpbxqdUTFccpH1Cw6YnV8lTWLyxJavbisombJCSqPc/jfSiur4wv/X0V1zNLS8qOtiiiJKVu17IiVUeWrjlW2qqC4bGVBydHKjzj8fA07/PfSeKoKikqrlheVxFN5jMKSqhWFJZXxFYdVFJ6gpKJwRfHRyguXFx1RuWrtnNpNmyeEbdzUdERdhuqjNh1jS8rqEmloTlt9Y2YajtFyos3paD2iKb7GDGxuajtiy7GaW7eNb2nd/gmzBwhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAACCkCcBAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAAEAQAgAAAAAAQBACAAAAAABAEAIAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAAQhAAAAAAAABCEAAAAAAAAEIQAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAAAAQQgAAAAAAABBCAAAAAAAAEEIAAAAAABAEPIkAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAAAIQgAAAAAAAAhCAAAAAAAACEIAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAAAAghAAAAAAAACCEAAAAAAAAIIQAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAAIAgBAAAAAAAgCAEAAAAAACAIAQAAAAAACEKeBAAAAAAAgHz2/1+2VRdzMnZPAAAAAElFTkSuQmCC"/>
  </defs>
 </g>
 <g transform="translate(0,2136)">
  <path d="m13 2.3213h0.8333c0.9167 0 1.6667 0.74731 1.6667 1.6607v11.625c0 0.9134-0.75 1.6607-1.6667 1.6607h-11.667c-0.925 0-1.6667-0.7473-1.6667-1.6607l0.008333-11.625c0-0.91338 0.73334-1.6607 1.6583-1.6607h0.83333v-1.6607h1.6667v1.6607h6.6666v-1.6607h1.6667v1.6607zm-10.833 13.285h11.667v-9.1338h-11.667v9.1338z" clip-rule="evenodd" fill="#5F6368" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,3506)" fill="#5F6368">
  <path d="m12.45 6.9344v-1.1791h1.175l3.5417-3.5207c-1.3-1.2953-3.0083-1.943-4.7167-1.943-1.7083 0-3.4083 0.64767-4.7166 1.943l-7.0667 7.0496v1.1708h1.175l3.5333-3.5207c0.975 0.97151 2.2583 1.4614 3.5333 1.4614 1.275 0 2.5666-0.4899 3.5416-1.4614zm-3.5333-3.529c0.94167-0.93829 2.2-1.4614 3.5333-1.4614 0.7584 0 1.4917 0.16607 2.1584 0.4816l-1.6667 1.6607h-2.1583v2.0676c-0.55 0.37366-1.1917 0.57294-1.8667 0.57294-0.89166 0-1.725-0.34874-2.3583-0.9715l2.3583-2.3499z"/>
  <path d="m15.667 12.116h-7.5c-0.45833 0-0.83333 0.3736-0.83333 0.8303v1.6607c0 0.4567 0.375 0.8303 0.83333 0.8303h7.5c0.4583 0 0.8333-0.3736 0.8333-0.8303v-1.6607c0-0.4567-0.375-0.8303-0.8333-0.8303z"/>
  <path d="m9.8337 9.6247c-0.45833 0-0.83333 0.37365-0.83333 0.83037v0.8303h5.8334v-0.8303c0-0.45672-0.375-0.83037-0.8334-0.83037h-4.1666z"/>
 </g>
 <g transform="translate(0,1792)">
  <path d="m12 4c-2.21 0-4 1.79-4 4s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm2 4c0-1.1-0.9-2-2-2s-2 0.9-2 2 0.9 2 2 2 2-0.9 2-2zm4 9c-0.2-0.71-3.3-2-6-2s-5.8 1.29-6 2.01v0.99h12v-1zm-14 0c0-2.66 5.33-4 8-4s8 1.34 8 4v3h-16v-3z" clip-rule="evenodd" fill="#5F6368" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,712)">
  <path d="m16.138 1.7963-1.2135-1.214c-0.7761-0.77636-2.0469-0.77636-2.8281 0l-11.37 11.374v4.0433h4.0417l11.37-11.374c0.7865-0.78157 0.7865-2.0529 0-2.8293zm-12.203 12.203h-1.2083v-1.2088l8.6614-8.665 1.2084 1.2088-8.6615 8.665zm4.7917 2.0008 4-4.0016h6v4.0016h-10z" fill="#174EA6"/>
 </g>
 <g transform="translate(0,1608)">
  <path d="m14.758 2.1917-1.95-1.9417c-0.325-0.325-0.8583-0.325-1.175 0l-1.1833 1.175-1.1833-1.175c-0.31667-0.325-0.85834-0.33333-1.1833-0.008333l-5.3083 5.3 1.1667 1.1667 4.7167-4.7167 0.60834 0.60833-2.1083 2.1083 3.1334 3.1333 4.475-4.4667c0.325-0.325 0.3166-0.85833-0.0084-1.1833zm-14.758 12.808v-3.125l6.275-6.275 3.125 3.125-6.2833 6.275h-3.1167z" clip-rule="evenodd" fill="#5F6368" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,2786)">
  <path d="m13.666 6.964-1.175-1.1708-4.6583 4.6334v-10.105h-1.6667v10.105l-4.65-4.6416-1.1833 1.1791 6.6667 6.6428 6.6666-6.6428z" fill="#174EA6"/>
 </g>
 <g transform="translate(0,3298)">
  <path d="M20 2H4c-1.1 0-1.99.9-1.99 2L2 22l4-4h14c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm-7 12h-2v-2h2v2zm0-4h-2V6h2v4z"/>
 </g>
 <g transform="translate(0,2160)">
  <defs>
   <filter id="drop-shadow">
    <feGaussianBlur in="SourceAlpha" stdDeviation="1.4"/>
    <feOffset dx="0" dy="1" result="offsetblur"/>
    <feFlood flood-color="rgba(0,0,0,0.8)"/>
    <feComposite in2="offsetblur" operator="in"/>
    <feMerge>
     <feMergeNode/>
     <feMergeNode in="SourceGraphic"/>
    </feMerge>
   </filter>
  </defs>
  <g fill="#fff" filter="url(#drop-shadow)">
   <rect x="3" y="8" width="4" height="4"/>
   <rect x="9" y="8" width="4" height="4"/>
   <rect x="15" y="8" width="4" height="4"/>
   <rect x="3" y="14" width="4" height="4"/>
   <rect x="9" y="14" width="4" height="4"/>
   <rect x="15" y="14" width="4" height="4"/>
  </g>
 </g>
 <g transform="translate(0,128)">
  <path d="M6 2c-1.1 0-1.99.9-1.99 2L4 20c0 1.1.89 2 1.99 2H18c1.1 0 2-.9 2-2V8l-6-6H6zm12 15.59l-2.2-2.2c.44-.69.7-1.51.7-2.39 0-2.48-2.02-4.5-4.5-4.5S7.5 10.52 7.5 13s2.02 4.5 4.5 4.5c.88 0 1.69-.26 2.39-.7l3.2 3.2H6V4h7.17L18 8.83v8.76zm-6-2.09a2.5 2.5 0 0 1 0-5 2.5 2.5 0 0 1 0 5z" fill="#fff"/>
 </g>
 <g transform="translate(0,1896)">
  <path d="M6 2c-1.1 0-1.99.9-1.99 2L4 20c0 1.1.89 2 1.99 2H18c1.1 0 2-.9 2-2V8l-6-6H6zm12 15.59l-2.2-2.2c.44-.69.7-1.51.7-2.39 0-2.48-2.02-4.5-4.5-4.5S7.5 10.52 7.5 13s2.02 4.5 4.5 4.5c.88 0 1.69-.26 2.39-.7l3.2 3.2H6V4h7.17L18 8.83v8.76zm-6-2.09a2.5 2.5 0 0 1 0-5 2.5 2.5 0 0 1 0 5z"/>
 </g>
 <g transform="translate(0,2930)">
  <path d="M12 17.27L18.18 21l-1.64-7.03L22 9.24l-7.19-.61L12 2 9.19 8.63 2 9.24l5.46 4.73L5.82 21z"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1672)">
  <path d="M12 17.27L18.18 21l-1.64-7.03L22 9.24l-7.19-.61L12 2 9.19 8.63 2 9.24l5.46 4.73L5.82 21z" fill="#fff"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,2016)">
  <path d="M20 2H4c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zM9 17c-2.8 0-5-2.2-5-5s2.2-5 5-5c1.3 0 2.4.5 3.3 1.3L11 9.6c-.3-.4-1-.8-2-.8-1.8 0-3.2 1.4-3.2 3.2s1.5 3.2 3.2 3.2c2 0 2.8-1.4 2.9-2.4H9V11h4.7c.06.29.1.7.1 1.1C13.8 15 11.9 17 9 17zm11-5h-2v2h-1v-2h-2v-1h2V9h1v2h2v1z" fill="#fff"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1368)">
  <path d="M20 2H4c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zM9 17c-2.8 0-5-2.2-5-5s2.2-5 5-5c1.3 0 2.4.5 3.3 1.3L11 9.6c-.3-.4-1-.8-2-.8-1.8 0-3.2 1.4-3.2 3.2s1.5 3.2 3.2 3.2c2 0 2.8-1.4 2.9-2.4H9V11h4.7c.06.29.1.7.1 1.1C13.8 15 11.9 17 9 17zm11-5h-2v2h-1v-2h-2v-1h2V9h1v2h2v1z"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,3138)">
  <g fill="#fff">
   <path d="m11 10c1.104 0 2-0.896 2-2s-0.896-2-2-2c-1.105 0-1.999 0.896-1.999 2s0.894 2 1.999 2zm0 1c-2 0-4 0.699-4 1.6v1.4h8v-1.4c0-0.901-2-1.6-4-1.6z"/>
   <circle cx="5.5" cy="9.5" r="1.5"/>
   <path d="m5.5 12.125c-1.25 0-2.5 0.437-2.5 1v0.875h5v-0.875c0-0.563-1.25-1-2.5-1z"/>
   <circle cx="16.5" cy="9.5" r="1.5"/>
   <path d="m16.5 12.125c-1.25 0-2.5 0.437-2.5 1v0.875h5v-0.875c0-0.563-1.25-1-2.5-1z"/>
  </g>
 </g>
 <g transform="translate(0,3058)">
  <path d="M4 4v2.01C5.83 3.58 8.73 2 12.01 2 17.53 2 22 6.48 22 12s-4.47 10-9.99 10C6.48 22 2 17.52 2 12h2c0 4.42 3.58 8 8 8s8-3.58 8-8-3.58-8-8-8C9.04 4 6.47 5.61 5.09 8H8v2H2V4h2z"/>
  <path d="M13 12V6h-2v7l4.97 3.49 1.26-1.55z"/>
 </g>
 <g transform="translate(0,448)">
  <path d="M10 4H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2h-8l-2-2z" fill="#FFF"/>
 </g>
 <g transform="translate(0,2722)">
  <path d="M13.6316 10C14.2311 10 14.7679 10.2829 15.0899 10.72L19 16L15.0899 21.28C14.7679 21.7171 14.2311 22 13.6316 22L3.78948 21.9914C2.80527 21.9914 2 21.2285 2 20.2857V11.7143C2 10.7714 2.80527 10.0086 3.78948 10.0086L13.6316 10ZM4 20H14L16.8078 16L14 12H8.5H4V20Z" clip-rule="evenodd" fill-rule="evenodd"/>
  <path d="m22.364 5.2727-0.5114-1.125-1.125-0.51138 1.125-0.51136 0.5114-1.125 0.5113 1.125 1.125 0.51136-1.125 0.51138-0.5113 1.125zm0 5.7273-0.5114-1.125-1.125-0.51136 1.125-0.51138 0.5114-1.125 0.5113 1.125 1.125 0.51138-1.125 0.51136-0.5113 1.125zm-4.091-1.2273-1.0227-2.25-2.25-1.0227 2.25-1.0227 1.0227-2.25 1.0228 2.25 2.2499 1.0227-2.2499 1.0227-1.0228 2.25zm0-1.9841 0.4091-0.87955 0.8796-0.4091-0.8796-0.40909-0.4091-0.87955-0.4091 0.87955-0.8795 0.40909 0.8795 0.4091 0.4091 0.87955z"/>
  <path d="m17.536 7.4818c0.5423 0 0.9819-0.43957 0.9819-0.98182 0-0.54224-0.4396-0.98182-0.9819-0.98182-0.5422 0-0.9818 0.43958-0.9818 0.98182 0 0.54225 0.4396 0.98182 0.9818 0.98182z"/>
  <path d="m19.991 6.5c0 0.54224-0.9305 0.98182-1.4727 0.98182-0.5423 0-0.9819-0.43958-0.9819-0.98182s-0.0513-1.4727 0.491-1.4727c0.5422 0 1.9636 0.9305 1.9636 1.4727z"/>
  <path d="m19.009 7.4817c0 0.27113-0.2198 0.49091-0.4909 0.49091s-0.4909-0.21978-0.4909-0.49091c0-0.27112 0.2198-0.49091 0.4909-0.49091s0.4909 0.21979 0.4909 0.49091z"/>
 </g>
 <g transform="translate(0,3034)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M17.63 5.84C17.27 5.33 16.67 5 16 5L5 5.01C3.9 5.01 3 5.9 3 7v10c0 1.1.9 1.99 2 1.99L16 19c.67 0 1.27-.33 1.63-.84L22 12l-4.37-6.16zM16 17H5V7h11l3.55 5L16 17z"/>
 </g>
 <g transform="translate(0,2970)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M17.63 5.84C17.27 5.33 16.67 5 16 5L5 5.01C3.9 5.01 3 5.9 3 7v10c0 1.1.9 1.99 2 1.99L16 19c.67 0 1.27-.33 1.63-.84L22 12l-4.37-6.16zM16 17H5V7h11l3.55 5L16 17z" fill="#fff"/>
 </g>
 <g transform="translate(0,2096)">
  <path d="M15.41 16.09l-4.58-4.59 4.58-4.59L14 5.5l-6 6 6 6z" fill="#fff"/>
  <path d="M0-.5h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,2264)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M3.9 12c0-1.71 1.39-3.1 3.1-3.1h4V7H7c-2.76 0-5 2.24-5 5s2.24 5 5 5h4v-1.9H7c-1.71 0-3.1-1.39-3.1-3.1zM8 13h8v-2H8v2zm9-6h-4v1.9h4c1.71 0 3.1 1.39 3.1 3.1s-1.39 3.1-3.1 3.1h-4V17h4c2.76 0 5-2.24 5-5s-2.24-5-5-5z"/>
 </g>
 <g transform="translate(0,472)">
  <path d="M18 8h-1V6c0-2.76-2.24-5-5-5S7 3.24 7 6v2H6c-1.1 0-2 .9-2 2v10c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V10c0-1.1-.9-2-2-2zM9 6c0-1.66 1.34-3 3-3s3 1.34 3 3v2H9V6zm9 14H6V10h12v10zm-6-3c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2z" fill="#fff"/>
 </g>
 <g transform="translate(0,3258)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M19 4H5c-1.11 0-2 .9-2 2v12c0 1.1.89 2 2 2h14c1.1 0 2-.9 2-2V6c0-1.1-.9-2-2-2zm-8 7H9.5v-.5h-2v3h2V13H11v1c0 .55-.45 1-1 1H7c-.55 0-1-.45-1-1v-4c0-.55.45-1 1-1h3c.55 0 1 .45 1 1v1zm7 0h-1.5v-.5h-2v3h2V13H18v1c0 .55-.45 1-1 1h-3c-.55 0-1-.45-1-1v-4c0-.55.45-1 1-1h3c.55 0 1 .45 1 1v1z" fill="#fff"/>
 </g>
 <g transform="translate(0,1856)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M19 4H5c-1.11 0-2 .9-2 2v12c0 1.1.89 2 2 2h14c1.1 0 2-.9 2-2V6c0-1.1-.9-2-2-2zm-8 7H9.5v-.5h-2v3h2V13H11v1c0 .55-.45 1-1 1H7c-.55 0-1-.45-1-1v-4c0-.55.45-1 1-1h3c.55 0 1 .45 1 1v1zm7 0h-1.5v-.5h-2v3h2V13H18v1c0 .55-.45 1-1 1h-3c-.55 0-1-.45-1-1v-4c0-.55.45-1 1-1h3c.55 0 1 .45 1 1v1z"/>
 </g>
 <g transform="translate(0,1936)">
  <path d="m7 10 5 5 5-5z" fill="#fff"/>
  <path d="M0 0h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,2746)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z" fill="#fff"/>
 </g>
 <g transform="translate(0,2056)">
  <path d="M4 15h16v-2H4v2zm0 4h16v-2H4v2zm0-8h16V9H4v2zm0-6v2h16V5H4z" fill="#fff"/>
 </g>
 <g transform="translate(0,1200)">
  <path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10zm-8.01-9l-1.41 1.41L12.16 12H8v2h4.16l-1.59 1.59L11.99 17 16 13.01 11.99 9z"/>
 </g>
 <g transform="translate(0,1568)">
  <path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10zm-8.01-9l-1.41 1.41L12.16 12H8v2h4.16l-1.59 1.59L11.99 17 16 13.01 11.99 9z" fill="#fff"/>
 </g>
 <g transform="translate(0,408)">
  <path d="m16.625 3.5h-12.25c-0.97125 0-1.75 0.7875-1.75 1.75v10.5c0 0.9625 0.77875 1.75 1.75 1.75h3.5v-1.75h-3.5v-8.75h12.25v8.75h-3.5v1.75h3.5c0.9625 0 1.75-0.7875 1.75-1.75v-10.5c0-0.9625-0.77875-1.75-1.75-1.75zm-6.125 5.25-3.5 3.5h2.625v5.25h1.75v-5.25h2.625l-3.5-3.5z" fill="#fff"/>
 </g>
 <g transform="translate(0,3530)">
  <path d="m16.625 3.5h-12.25c-0.97125 0-1.75 0.7875-1.75 1.75v10.5c0 0.9625 0.77875 1.75 1.75 1.75h3.5v-1.75h-3.5v-8.75h12.25v8.75h-3.5v1.75h3.5c0.9625 0 1.75-0.7875 1.75-1.75v-10.5c0-0.9625-0.77875-1.75-1.75-1.75zm-6.125 5.25-3.5 3.5h2.625v5.25h1.75v-5.25h2.625l-3.5-3.5z"/>
 </g>
 <g transform="translate(0,1328)">
  <path d="m22.051 12.838v-4.755c0-4.464-3.619-8.083-8.083-8.083s-8.083 3.619-8.083 8.083v4.754c-0.678 0.106-1.201 0.695-1.201 1.401v12.342c0 0.781 0.639 1.42 1.42 1.42h15.72c0.781 0 1.42-0.639 1.42-1.42v-12.342c0-0.703-0.519-1.29-1.193-1.4zm-8.083-9.561c2.594 0 4.697 2.103 4.697 4.697v4.844h-9.394v-4.844c0-2.594 2.103-4.697 4.697-4.697zm1.093 17.549v3.642h-2.258v-3.7c-0.717-0.412-1.201-1.185-1.201-2.07 0-1.317 1.068-2.385 2.385-2.385s2.385 1.067 2.385 2.385c-1e-3 0.929-0.534 1.736-1.311 2.128z" fill="#aaa"/>
 </g>
 <g transform="translate(0,368)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M19 19H5V5h7V3H5c-1.11 0-2 .9-2 2v14c0 1.1.89 2 2 2h14c1.1 0 2-.9 2-2v-7h-2v7zM14 3v2h3.59l-9.83 9.83 1.41 1.41L19 6.41V10h2V3h-7z"/>
 </g>
 <g transform="translate(0,2304)">
  <path d="M0 0h24v24H0z" fill="none"/>
  <path d="M19 19H5V5h7V3H5c-1.11 0-2 .9-2 2v14c0 1.1.89 2 2 2h14c1.1 0 2-.9 2-2v-7h-2v7zM14 3v2h3.59l-9.83 9.83 1.41 1.41L19 6.41V10h2V3h-7z" fill="#fff"/>
 </g>
 <g transform="translate(0,3426)">
  <path d="M19 8h-1V3H6v5H5c-1.66 0-3 1.34-3 3v6h4v4h12v-4h4v-6c0-1.66-1.34-3-3-3zm-3 11H8v-4h8v4zm0-11H8V5h8v3zm2 4.5c-.55 0-1-.45-1-1s.45-1 1-1 1 .45 1 1-.45 1-1 1z" fill="#fff"/>
 </g>
 <g transform="translate(0,512)">
  <path d="M19 8h-1V3H6v5H5c-1.66 0-3 1.34-3 3v6h4v4h12v-4h4v-6c0-1.66-1.34-3-3-3zm-3 11H8v-4h8v4zm0-11H8V5h8v3zm2 4.5c-.55 0-1-.45-1-1s.45-1 1-1 1 .45 1 1-.45 1-1 1z"/>
 </g>
 <g transform="translate(0,168)">
  <path d="m10.5 3.5c-3.59 0-6.5 2.91-6.5 6.5s2.91 6.5 6.5 6.5 6.5-2.91 6.5-6.5-2.91-6.5-6.5-6.5zm3.303 8.937h-1.678v-0.812s0-1.625-1.625-1.625h-2.438l0.01-1.625h0.789c0.543 0 0.826 0 0.826-0.711v-0.914h0.865c1.572 0 1.572-1.625 1.572-1.625v-0.38c2.241 0.695 3.875 2.787 3.875 5.255 0 1.423-0.548 2.717-1.438 3.694v-0.478c1e-3 -0.556-0.203-0.779-0.758-0.779zm-8.803-2.437c0-0.73 0.146-1.427 0.405-2.064l1.032 2.064s3.25 2.43 3.25 2.438v0.742c0 0.883 0.812 0.811 0.812 0.883v1.438c-3.031-1e-3 -5.499-2.468-5.499-5.501z" fill="#fff"/>
 </g>
 <g transform="translate(0,976)">
  <path d="m18.41 5.8-1.21-1.21c-0.78-0.78-2.05-0.78-2.83 0l-11.37 11.37v4.04h4.04l11.37-11.37c0.79-0.78 0.79-2.05 0-2.83zm-12.2 12.2h-1.21v-1.21l8.66-8.66 1.21 1.21-8.66 8.66zm4.79 2 4-4h6v4h-10z"/>
 </g>
 <g transform="translate(0,856)">
  <path d="m18.41 5.8-1.21-1.21c-0.78-0.78-2.05-0.78-2.83 0l-11.37 11.37v4.04h4.04l11.37-11.37c0.79-0.78 0.79-2.05 0-2.83zm-12.2 12.2h-1.21v-1.21l8.66-8.66 1.21 1.21-8.66 8.66zm4.79 2 4-4h6v4h-10z" fill="#fff"/>
 </g>
 <g transform="translate(0,3098)">
  <path d="M15.73 3H8.27L3 8.27v7.46L8.27 21h7.46L21 15.73V8.27L15.73 3zM19 14.9L14.9 19H9.1L5 14.9V9.1L9.1 5h5.8L19 9.1v5.8z"/>
  <circle cx="12" cy="16" r="1"/>
  <path d="m11 7h2v7h-2z"/>
 </g>
 <g transform="translate(0,3714)" fill="#fff">
  <path d="M15.73 3H8.27L3 8.27v7.46L8.27 21h7.46L21 15.73V8.27L15.73 3zM19 14.9L14.9 19H9.1L5 14.9V9.1L9.1 5h5.8L19 9.1v5.8z"/>
  <circle cx="12" cy="16" r="1"/>
  <path d="m11 7h2v7h-2z"/>
 </g>
 <g transform="translate(0,2504)">
  <g fill-rule="evenodd" xmlns:sketch="http://www.bohemiancoding.com/sketch/ns">
   <path d="m2.0044 6.6876 1.2789 2.2832 9.5747-8.9708 1.142 2.2593-10.218 9.7407-3.782-3.9102 2.0044-1.4022z" fill="#c1bfbf"/>
  </g>
 </g>
 <g transform="translate(0,3594)">
  <path d="M4 4v2.01C5.83 3.58 8.73 2 12.01 2 17.53 2 22 6.48 22 12s-4.47 10-9.99 10C6.48 22 2 17.52 2 12h2c0 4.42 3.58 8 8 8s8-3.58 8-8-3.58-8-8-8C9.04 4 6.47 5.61 5.09 8H8v2H2V4h2zm9 8V6h-2v7l4.97 3.49 1.26-1.55L13 12z" clip-rule="evenodd" fill="#fff" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,248)">
  <path d="M8.59 16.34l4.58-4.59-4.58-4.59L10 5.75l6 6-6 6z" fill="#fff"/>
  <path d="M0-.25h24v24H0z" fill="none"/>
 </g>
 <g transform="translate(0,1752)">
  <polygon points="11 14 4.5 7.5 6 6 11 11 16 6 17.5 7.5" fill="#fff"/>
 </g>
 <g transform="translate(0,3754)">
  <polygon points="11 6 4.5 12.5 6 14 11 9 16 14 17.5 12.5" fill="#fff"/>
 </g>
 <g transform="translate(0,2682)">
  <g transform="matrix(.69989 0 0 .69989 -.91859 3.0615)" fill="#fff">
   <path d="m19.802 30.409-5.5907-5.5907-1.8971 1.8971 7.4878 7.4878 16.088-16.088-1.8971-1.8971-14.191 14.191z" fill="#fff"/>
  </g>
 </g>
 <g transform="translate(0,592)">
  <path d="M13.85 22.25h-3.7c-.74 0-1.36-.54-1.45-1.27l-.27-1.89c-.27-.14-.53-.29-.79-.46l-1.8.72c-.7.26-1.47-.03-1.81-.65L2.2 15.53c-.35-.66-.2-1.44.36-1.88l1.53-1.19c-.01-.15-.02-.3-.02-.46 0-.15.01-.31.02-.46l-1.52-1.19c-.59-.45-.74-1.26-.37-1.88l1.85-3.19c.34-.62 1.11-.9 1.79-.63l1.81.73c.26-.17.52-.32.78-.46l.27-1.91c.09-.7.71-1.25 1.44-1.25h3.7c.74 0 1.36.54 1.45 1.27l.27 1.89c.27.14.53.29.79.46l1.8-.72c.71-.26 1.48.03 1.82.65l1.84 3.18c.36.66.2 1.44-.36 1.88l-1.52 1.19c.01.15.02.3.02.46s-.01.31-.02.46l1.52 1.19c.56.45.72 1.23.37 1.86l-1.86 3.22c-.34.62-1.11.9-1.8.63l-1.8-.72c-.26.17-.52.32-.78.46l-.27 1.91c-.1.68-.72 1.22-1.46 1.22zm-3.23-2h2.76l.37-2.55.53-.22c.44-.18.88-.44 1.34-.78l.45-.34 2.38.96 1.38-2.4-2.03-1.58.07-.56c.03-.26.06-.51.06-.78s-.03-.53-.06-.78l-.07-.56 2.03-1.58-1.39-2.4-2.39.96-.45-.35c-.42-.32-.87-.58-1.33-.77l-.52-.22-.37-2.55h-2.76l-.37 2.55-.53.21c-.44.19-.88.44-1.34.79l-.45.33-2.38-.95-1.39 2.39 2.03 1.58-.07.56a7 7 0 0 0-.06.79c0 .26.02.53.06.78l.07.56-2.03 1.58 1.38 2.4 2.39-.96.45.35c.43.33.86.58 1.33.77l.53.22.38 2.55z"/>
  <circle cx="12" cy="12" r="3.5"/>
 </g>
 <g transform="translate(0,3218)">
  <path d="M9 12c2.21 0 4-1.79 4-4s-1.79-4-4-4-4 1.79-4 4 1.79 4 4 4zm0-6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2zm0 7c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4zm6 5H3v-.99C3.2 16.29 6.3 15 9 15s5.8 1.29 6 2v1zm3-4v-3h-3V9h3V6h2v3h3v2h-3v3h-2z" fill="#fff"/>
 </g>
 <g transform="translate(0,2994)">
  <path d="M9 12c2.21 0 4-1.79 4-4s-1.79-4-4-4-4 1.79-4 4 1.79 4 4 4zm0-6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2zm0 7c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4zm6 5H3v-.99C3.2 16.29 6.3 15 9 15s5.8 1.29 6 2v1zm3-4v-3h-3V9h3V6h2v3h3v2h-3v3h-2z"/>
 </g>
 <g transform="translate(0,3674)">
  <metadata id="metadata19" xmlns:cc="http://creativecommons.org/ns#" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
   <rdf:RDF>
    <cc:Work rdf:about="">
     <dc:format>image/svg+xml</dc:format>
     <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
    </cc:Work>
   </rdf:RDF>
  </metadata>
  <!-- Generator: Sketch 39.1 (31720) - http://www.bohemiancoding.com/sketch -->
  <title id="title4">ic_my_drive_black_48dp copy</title>
  <desc id="desc6">Created with Sketch.</desc>
  <g id="ASSETS" transform="matrix(.3125 0 0 .3125 .0021186 .070829)" fill="none">
   <g id="icons" transform="translate(-275,-4)">
    <g id="ic_my_drive_black_48dp-copy" transform="translate(269)">
     <g id="Group">
      <path id="Shape" d="m0 0h48v48h-48v-48zh48v48h-48v-48z"/>
      <path id="path15" d="m6 40.02c0 2.2 1.79 3.98 3.99 3.98h28.02c2.2 0 3.99-1.8 3.99-3.98v-4.02h-36v4.02zm30-2.02c1.1 0 2 0.9 2 2s-0.9 2-2 2-2-0.9-2-2 0.9-2 2-2zm2.01-34h-28.02c-2.2 0-3.99 1.8-3.99 3.98v26.02h36v-26.02c0-2.2-1.79-3.98-3.99-3.98z" fill="#8f8f8f"/>
     </g>
    </g>
   </g>
  </g>
 </g>
 <g transform="translate(0,64)">
  <path d="m23 21-11-19-11 19h22zm-12-3v-2h2v2h-2zm0-4h2v-4h-2v4z" clip-rule="evenodd" fill="#F9AB00" fill-rule="evenodd"/>
 </g>
 <g transform="translate(0,776)">
  <path d="M15.5 14h-.79l-.28-.27C15.41 12.59 16 11.11 16 9.5 16 5.91 13.09 3 9.5 3S3 5.91 3 9.5 5.91 16 9.5 16c1.61 0 3.09-.59 4.23-1.57l.27.28v.79l5 4.99L20.49 19l-4.99-5zm-6 0C7.01 14 5 11.99 5 9.5S7.01 5 9.5 5 14 7.01 14 9.5 11.99 14 9.5 14z" fill="#fff"/>
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M12 10h-2v2H9v-2H7V9h2V7h1v2h2v1z" fill="#fff"/>
 </g>
 <g transform="translate(0,2200)">
  <path d="M19 13H5v-2h14v2z" fill="#fff"/>
 </g>
 <g transform="translate(0,1016)">
  <path d="M0 0h24v24H0V0z" fill="none"/>
  <path d="M15.5 14h-.79l-.28-.27C15.41 12.59 16 11.11 16 9.5 16 5.91 13.09 3 9.5 3S3 5.91 3 9.5 5.91 16 9.5 16c1.61 0 3.09-.59 4.23-1.57l.27.28v.79l5 4.99L20.49 19l-4.99-5zm-6 0C7.01 14 5 11.99 5 9.5S7.01 5 9.5 5 14 7.01 14 9.5 11.99 14 9.5 14zM7 9h5v1H7z" fill="#fff"/>
 </g>
 <g transform="translate(0,552)">
  <path d="M19 13h-6v6h-2v-6H5v-2h6V5h2v6h6v2z" fill="#fff"/>
 </g>
</svg>

------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/css
Content-Transfer-Encoding: binary
Content-Location: https://www.gstatic.com/og/_/ss/k=og.qtm.Bcf36HdLxAc.L.W.O/m=qcwid/excm=qaaw,qadd,qaid,qein,qhaw,qhba,qhbr,qhch,qhga,qhid,qhin/d=1/ed=1/ct=zgms/rs=AA2YrTtrdJEPAVAbPPca5uf3TCfVu9JrgA

@charset "utf-8";

.gb_4e { background: rgba(60, 64, 67, 0.9); border-radius: 4px; color: rgb(255, 255, 255); font: 500 12px / 16px Roboto, arial, sans-serif; letter-spacing: 0.8px; margin-top: 4px; min-height: 14px; padding: 4px 8px; position: absolute; z-index: 1000; -webkit-font-smoothing: antialiased; }

.gb_Ic { text-align: left; }

.gb_Ic > * { color: rgb(189, 193, 198); line-height: 16px; }

.gb_Ic div:first-child { color: white; }

sentinel { }
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/jpeg
Content-Transfer-Encoding: binary
Content-Location: https://lh3.googleusercontent.com/ogw/AOLn63Fd7vZE5o2FaKK7Sg0PDYjfXo_g8YLZTYOwvcVc=s32-c-mo

���� JFIF      �� ~Exif  II*     1    &   i�    .       Google    �    0220�       �    X             R98      0100    �� � 


		��  @ @ ��             	�� 0      ! 1"AQaq2��#�b����                 ��                 ��   ? ��6�[Ԛ|Y,�r��BV�ҽ�(c�@����J�
#mš)Jp[���A����(�]��K�(C�'�?���O_ظe?��;zi8bD����3�<{���O5�_�m��JU��	���zQjv�x#<���A:ϯT.�:��k��Ni��	KNv��@� ���=ڶ�&�H�R很��N0���6�{	e=�0�/zBR�NV8� �oQ���Qݭ&E-�e�Q�Cn��AB�p���5ѯ����ڈ����n���).gbF  ����M������%�:2JO>��U�y��=خ-���� ��� ��N��%KRZPK	8H'�9���՛1s)N�U(��T�>�.p�R�� }� ��nh!� �iiǦ9NafrX�)�ê[�pq[T�T
Rd��z�����D��M��n�N�4�џo�Y'�78J�y��>�����L���-���c�?T��vP�m�
o|����%(
'%I ���t�^�N�W%t:��]�Хび �O���>\z����3�$�ˏ(c�
�?*�ǲGA��f"�,4���h4�o@;�������v�ܠ�6�@Y�>��AM}�:R����Jn#��%��>�:�C�NgԒ���G�@�ڻh�D3m��܌Ȗ�o0���o)qCjЕ�g��c��c�5�I��L�3��)tvX�*��]�Tҵ���JNJ]J��<��`��z
�T�V^�p�_�U��n�Gra����Ys���%��6�%CjE;Ln�=�����-������Ф*:r�
�#i�$a�A�z��_�*�NnAu�-=�YaǊ��Vԅ(ダ9�ӂ������mE�<��-�-�[�x<��@� )_��5���(��B��	S-zB�?n|s�i���n�������k[Ҟ��%Ѵ�w�pT@>=��{�n��V�i�d&jWO�E�8)�"J�+� �ڷ)���p�����������1��N�ó#�y	i/I���hF0�)�7��W ��m�A�B5�7�X����P_�!O:�p�w8N��}�=N�B���0hKJ�>��-�'�����ܯ�$���
ХX_���z�2�J�R�ox���O���O�<x�-5cB)7]U$��Q)��l�H�����	P�pp	�1���'m7^j;�
�-ID�ܪ�A��ʚgi�/
9Io�$�bЁjȩ*֥R�H�T_}m[�P�' H���A{�iM�m*R���c�BВ���'$���=Ŷ�ȑ*[���R�D�׹Y[�������Ax)1݀aͪ)�T�$��C�~�O�}:v?���*
nZ�h����En�{
wԼo@�y�e	뜌 ���� ���mV�"�S��o�^T[J�� �9���jY�T�K�VA�Ug(1�G���㜏�Z��u߶h�(L�c��vz䥵=(�܇;��'{${c#'"������)�����.!����B�J�I��q��;�z���Zy�]�9������w!
N����� �:��|P��n�Bxʉ�q���-�˨8R��O��!I ��z=[�x�S6�Nj��b�Pu���%���R��8IQ� ���s��|�N�06����t�,j�$@�5�{2��H���m嬡���� z
IM�-�^�O�*�$+k�Jh��PFS��;|dx?N�G[��gW�a]��c���/b�S�;q�#?���|OjQj�����ڍ1P�ڔ6�q���������R��,��?c���6����.���Ҹ̘�S���_y
Q�$����AU�N��պ���\xJD,�@�
��-J�2�>��v�I���q-�탞�=2{����C�[�$�iݐ���$��A�uN�R��zDZv��i�Ө�S�@9a�:��Ϥ)**P�@�F��W���Z��?q��F{xhgQ��8󌎀Pڔd� #ߠ��O'����Ƈ��mD���T��u�0JgzA?A�_�U�T&ɇBL���*������u{���?��
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/png
Content-Transfer-Encoding: binary
Content-Location: https://drive-thirdparty.googleusercontent.com/32/type/application/x-virtualbox-vhd

�PNG

   IHDR           szz�    cHRM  z%  ��  ��  ��  u0  �`  :�  o�_�F   tIDATW�α�0DQ��,���8���.B�\gQ�����E��M�/[�s��}����(�(�Q�"� A�)�'D��H�!�W��,�P �  � �
p ��=X��Y    IEND�B`�
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/jpeg
Content-Transfer-Encoding: binary
Content-Location: https://lh3.googleusercontent.com/a/AAcHTtdQDe6r_XGCNEiOx6KZzpjviLw9RqZeAy_GGnpv=s50-c-k-no

���� JFIF      �� ~Exif  II*     1    &   i�    .       Google    �    0220�       �    X             R98      0100    �� � 


		��  2 2 ��              	�� 5       !1"Aq2a�#Q��B��$5RS��                 ��                 ��   ? �[
׶iU:[
S2d9�}�� �`���"��|S\����yԃ�� �����R���ՋZ�y��v���X_�Nכ�b��B�� �Oq�"�r�n�~Mj˫QnH����C.Gu���+�0�>��F�N]ӪW�(Q���챏.ؾ%Id$t��H�s�q�o뎿�N]^�Nj���Zqk��4�7,�_R	H��Gĕ6$�Xv�X6���� A����h&�W�{��T*US��Lw��� � |�sq��(�����W�^�Bn`e譇��ܐzg��8#x�	J���� �Na^�m ��d_<2�RQ9�t��*,�+;T�D�	냌��o@tK��TfDuչ���1��4�����P�T�E=IQRA�r2�N�p[R����&ڪ���3��b�2���8�)-�h2�6m)J�>e��y�l_��������:���6�nm\��:�h%k2j���d����c�(6P��k4����nP�lu�pO���ʬ]3�9��͗�u�$����l}p ޷��kwE3C�2B�7���:	�J����
%jW���qqi˘�<��oqIJ�y�{���d�T[�C���l�%�ϔ4��i���j (�m$~�נ���R6Dj�kU�TU��UG����R���S�)=
GQ�Q&�y�[�*0[_�1^��Kd�Q2�$v'�r�ε/v��ėH�jl��.:ۮ��S�Kd��?#����Ɓ]�X���P<9��6lw���x��u\����������D�])D����&��l����
8�׻(AQ�@Ϩ�;�{û~�f���Q��h�Yq��j|ͤж~`	?���R#�gb�	�|��������K��$`�#�΂F޷i�i�M��-��pW��8?�������o��\����)E�Ԟ羃4��C�T�&]FK��_���IPq����ԓ�،�8I���	*���%�UA�H�;х$�>�z��t�v���o*�k2)��i���R26��Nq�+9��q�S�|�l~�U�Ub"�y���椷�������#>�,�:�B�:�65Mh�C�8y����%!a=�A
8���q^�6�U�CJ��Kp9�(S����H�����C5���W&���n� j���נ��})��ڏ�sJ�}�3�5�i�+ƘiU��A�Rc
�����an%.�PFV���NjJNJ
�v��V��S$Z�g�`�ߋm;R�2v�$�$�@=z�;߈5��_�Ŗ#��JH��M ���q�1��}4�VLKFɵ��B�������s�~�˳K�J&2�@�AW�� ��=9�n��|yx�����mC�
^�3���▝�m�̰�L
)m��N��z��h3�i%���9m�i%@RAצ�H8�[ći7�.u��?a��[G�wʟ��}t��
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/png
Content-Transfer-Encoding: binary
Content-Location: https://drive-thirdparty.googleusercontent.com/16/type/application/vnd.google-apps.folder+shared

�PNG

   IHDR         ��a   gAMA  ���a   �IDAT8c`h�r��	������c��Å�@,�AR���� . vP�\
��o���<��Iy�$�2��������D��H����������h����w�ԩSy@4�,����Xj���W+69b�0���IMZZ�D��lA�ͷ���&�\�!��`:`�ya+�Dhr��`<�J�m7͘z
-    IEND�B`�
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: image/jpeg
Content-Transfer-Encoding: binary
Content-Location: https://lh3.googleusercontent.com/a/AAcHTtdQDe6r_XGCNEiOx6KZzpjviLw9RqZeAy_GGnpv=s64

���� JFIF      �� ~Exif  II*     1    &   i�    .       Google    �    0220�       �    X             R98      0100    �� � 


		��  @ @ ��             	�� 0      ! 1"AQaq2��#�b����                 ��                 ��   ? ��6�[Ԛ|Y,�r��BV�ҽ�(c�@����J�
#mš)Jp[���A����(�]��K�(C�'�?���O_ظe?��;zi8bD����3�<{���O5�_�m��JU��	���zQjv�x#<���A:ϯT.�:��k��Ni��	KNv��@� ���=ڶ�&�H�R很��N0���6�{	e=�0�/zBR�NV8� �oQ���Qݭ&E-�e�Q�Cn��AB�p���5ѯ����ڈ����n���).gbF  ����M������%�:2JO>��U�y��=خ-���� ��� ��N��%KRZPK	8H'�9���՛1s)N�U(��T�>�.p�R�� }� ��nh!� �iiǦ9NafrX�)�ê[�pq[T�T
Rd��z�����D��M��n�N�4�џo�Y'�78J�y��>�����L���-���c�?T��vP�m�
o|����%(
'%I ���t�^�N�W%t:��]�Хび �O���>\z����3�$�ˏ(c�
�?*�ǲGA��f"�,4���h4�o@;�������v�ܠ�6�@Y�>��AM}�:R����Jn#��%��>�:�C�NgԒ���G�@�ڻh�D3m��܌Ȗ�o0���o)qCjЕ�g��c��c�5�I��L�3��)tvX�*��]�Tҵ���JNJ]J��<��`��z
�T�V^�p�_�U��n�Gra����Ys���%��6�%CjE;Ln�=�����-������Ф*:r�
�#i�$a�A�z��_�*�NnAu�-=�YaǊ��Vԅ(ダ9�ӂ������mE�<��-�-�[�x<��@� )_��5���(��B��	S-zB�?n|s�i���n�������k[Ҟ��%Ѵ�w�pT@>=��{�n��V�i�d&jWO�E�8)�"J�+� �ڷ)���p�����������1��N�ó#�y	i/I���hF0�)�7��W ��m�A�B5�7�X����P_�!O:�p�w8N��}�=N�B���0hKJ�>��-�'�����ܯ�$���
ХX_���z�2�J�R�ox���O���O�<x�-5cB)7]U$��Q)��l�H�����	P�pp	�1���'m7^j;�
�-ID�ܪ�A��ʚgi�/
9Io�$�bЁjȩ*֥R�H�T_}m[�P�' H���A{�iM�m*R���c�BВ���'$���=Ŷ�ȑ*[���R�D�׹Y[�������Ax)1݀aͪ)�T�$��C�~�O�}:v?���*
nZ�h����En�{
wԼo@�y�e	뜌 ���� ���mV�"�S��o�^T[J�� �9���jY�T�K�VA�Ug(1�G���㜏�Z��u߶h�(L�c��vz䥵=(�܇;��'{${c#'"������)�����.!����B�J�I��q��;�z���Zy�]�9������w!
N����� �:��|P��n�Bxʉ�q���-�˨8R��O��!I ��z=[�x�S6�Nj��b�Pu���%���R��8IQ� ���s��|�N�06����t�,j�$@�5�{2��H���m嬡���� z
IM�-�^�O�*�$+k�Jh��PFS��;|dx?N�G[��gW�a]��c���/b�S�;q�#?���|OjQj�����ڍ1P�ڔ6�q���������R��,��?c���6����.���Ҹ̘�S���_y
Q�$����AU�N��պ���\xJD,�@�
��-J�2�>��v�I���q-�탞�=2{����C�[�$�iݐ���$��A�uN�R��zDZv��i�Ө�S�@9a�:��Ϥ)**P�@�F��W���Z��?q��F{xhgQ��8󌎀Pڔd� #ߠ��O'����Ƈ��mD���T��u�0JgzA?A�_�U�T&ɇBL���*������u{���?��
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic----
Content-Type: text/html
Content-ID: <frame-8DF312FC58F6EE99A3ED96B5411FF620@mhtml.blink>
Content-Transfer-Encoding: binary
Content-Location: https://clients6.google.com/static/proxy.html?usegapi=1&jsh=m%3B%2F_%2Fscs%2Fabc-static%2F_%2Fjs%2Fk%3Dgapi.gapi.en.K1LWthAzeb4.O%2Fd%3D1%2Frs%3DAHpOoo-TQTqnv7hwijrseP4JKJ1XY83Ehg%2Fm%3D__features__#parent=https%3A%2F%2Fdrive.google.com&rpctoken=361754389

<!DOCTYPE html><html><head><meta http-equiv="Content-Type" content="text/html; charset=windows-1252">
<title></title>
<meta http-equiv="X-UA-Compatible" content="IE=edge">


</head>
<body>


</body></html>
------MultipartBoundary--4O9EdP8RxyRaVerzT9q3vsReS9sglFW99GICny7Yic------
